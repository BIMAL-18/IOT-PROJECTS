PK   !l�Y^!H��  �a     cirkitFile.json�\[o�6�+���X.m/�=��'�t���$��ֱ��r.{���$}�/��d�5�����o>G��f��h������VM��.1�dw��>��V4ɖ�bַ�_;���.���y�ei�_���gu����K+dΪ��R*�eiM�K�������v�juS'0u
Sg0uS0u	SW0u�v@�a �Gސ�-l�)*r�-��,WVWym3�F��~�!C���Mō�T�Z�nh�L����X�qe,E��x�D<�U����Q�&�iK���6�q�q�q=[�1N��/mx��	C���DC"vl�H��c��!C�C)�� CK���Q�>�Q��1�	@�m�x�0PdhPdhP�b$�0�����W�����oPx�'���VH+4���
ObE$�"�XQI��4�K�4��i��~��r4ra��f��3i���@���am��y��8�I�D��$�44LҠ��!b���I@��QHL�5�-+�H]%����
~�&b� �Y"�:q~�bo	�<���;���%��pv�����)6�?���||����z՛�BS�}�;3��p+$���
Kb�'�"�X�I��$Vt�%o��4��i��� �A0Na��8�q�4(&�88�I�4(&iPLҠ��A1I�b�,��Sk��g1�Zí<����n�Y�F��g�D��p+��ttj����.�^����f=k��٥�d��ήf˹)m5s�w�U��.�A�yH��N@�yHlA�vd�Ь)(r@C3P����\\�>�菒����٬a����-�t������,�!�vN�����a I������x d� 	��Cb,O �]���	bH�o����9MW=4�]Ut����lW2}h*h�t,�B�	P��P��P_�P_C� �
�P�D����0��ydo�`�/z�&(N�<�7�3� 
� ��b�Q(�	�I	�J	�J�ʦ��y�l�f�y�]�LhG�Bt�3��+�#�]�蟁st}3�X�.t�A3��ydr���(E�@O��8ɞ�4�Ϟ���O�c������1��o���_E������x��8�^{�p5�S��� \԰W�^�xl{�5�� ^�x�5��f�U��w�_2"��Ԉ�8��z	��+8[�d�������d�c󐯡�1��SƇ}IV�>�4ؗ0`U�S
�}9V?�gطD@E������)���i�g?�����iȄ.|�E6]䴋n��i�t��.�����|>+:k��5�/4��lެ�5E���i���k����vi������VkWM~
��I<TRL��a9��J�,�5W9�TYS�U�[]�Jf�$4�L��"m��k����oL2w6�fQ�E�P���gŬ����vӕs���5d�|U��k*�i�%�6h�܊0$����d���(��܍��&z� dh@t�����j���D'[Q�Àniw-d-��y)�vDν�X���׶]�q%��ng��MSQ6�M�tҍ��,��G���`@*:����1����d��R�y�W�\HoG��ڐCꈀ
�2:�ۣ�EhݦŰ��97�x��xO\�~�D�8�w��p��<u�3��㷦��?TM���O�:&y6����R��D�ԃZ���>�Z��F27�B92u�+Q�܉I���&��r�:Lz:�>���|;���4�k�B!�tVL��qVL��5�G��+���A1�����X�����9����W��|�����d�7��7ۗw7��&k��RaR:�f��n��67��HMk��~�����l���~�n�+�ꂛ�5r�
�F�*We������A׏��G�r�c�+]�����
n�+�
ɍRX���-������]yi�v�|n��s漕؝�z�p�z����&~rk�tk3_ٽ�|�̫=˴*���#�pG�q琪�:1�=���`)�7]���v�gE+�c�R�JU�l��²�5�4.%+)V���+�RTذ��-��.�(r�"ՅfEA�
o����YT޹˾{�S�<J��g�o���~��[X��\�]�����j��{���g����4M���jw��/�P9SZ�!$G�U����C��pCs���e�mn-x��3�˺BhQ����?˹�х�&'�k'�`.�G����Ee��1�\W��$��BYU�ԜGT�~{�}l��be���_�z���fqq��n��/�C����w����������K'��{\���v�νif:������˾����ܖ�#�4��l�O��^��|��;e���ɢ�2G�MSG7����iR�p�1w[j�*��ܺ GRG%Q���D1�Y��ñ�����o�N*w/�Φ!�RJt�m�s�����aQ��M�.]�d�~;���}fS)���OM�߹6���EZ(�����;/��[aF��j>R�r`�אLyg��v�������_�����.����C��n����2gnٻ��Yl"���5?,���"%�Vg>}H雳�cB��m��L��������}}�;>�]��u�[/���U���T۷^`2$�2���N�g�/��j�w������-�R�ĕoF�}t���& fq����|{[�&̳Äs���R�q�@�%=�X�	@�R��Q
�r�?;��_&Lɲ4!�eb��i�/_ŲJư��/��\j@�R�K�~��=x�������a�a�e��F���8�<D^.�g����R���?щᏒ���K��!��q$�٠Q��"z��0{���S��%R��]��BJȊ��MCV�el���j��	���},5��Aj�QR\���F
����x��i&>r�?ґ2�My�c�s��W9��\�岃�x$5�yZ�Bj���.|�RxP���g�T,d׿N��)����*�2�C)"�7��QRc���C�H��������Lo���W٥G�*�i�g�����̿k�����?�����\v�l��`We�,7U����PK   lg�YG���F"  A"  /   images/07631829-c1ba-46e6-b58f-b7cc9d810cbd.pngA"�݉PNG

   IHDR   d   J   MD�   	pHYs  �v  �vU��   tEXtSoftware www.inkscape.org��<  !�IDATx��]y��U�?_��d�-�̄d�@  �(h�E���k�+RV)���O�R�JD|��|  !H� 	BL�>�Ifߺg�齧��w~�����2Y��y+]��}߹�~g?�{c!��N9��h���ifs�

���#-��0o;�z���@q~�Y�ߊ��nw�K[hv6�/��6zxn���e~��rMO�E�Qz�[�@����XL�C?)�f�a�;Q*++�;�x3�x�*-������W����_�=��I��L�O�%}��e�|yCl>z�0�0��[ISSgJ=��l5C�V����|�-��7���j�'��?�KO=�E�P��N%%�c�-t���uuŴeˍt����o��+fz��]_ob���������FFF�������	�����'�Uz25 ���"Z���B�p�FG�cO�3D21s�xC�-Bk����O��Y���PBo{+�r˃��?�L��@�0�v�R��ܾ�7�����_�ד(��N�BPE�������;��	�FΈ@��?��>��V����e	|���ut��#]xa%K�jVC*/���P?=�� =��|R?K��b$���~���M��^Q�[A0{+�p��Ӿ�UL�>z��8���&����f�9�����Yr�81ή�YN1r;�.�����?_���5|8�Y��SS����|41�Ç��t���R6#�ڤ�����ח���D�=�AyBb|
�9�]Rb�׳瓓QFZ�	��i���i#y���Ue)ӹoi&r:�X�{��9<�b�V�ҋ�a!�-7��(Uͩ�F�;ѱcc,��Y;;xp��B3��?��0΋�v�,�C��	��-�|�����R���Y�#U� ���t�@�`C4��_������B*80B=t�������Ɣ�i�u����"t�T�5Uc H?��t�}�2>���a�wR&���f������/��׳J(��y�~6z�n=����\����DA��
�����y&H8o��
8
ѨI����$���hٲ������x�b�z��Y.����iϞ1NUU��2��w� O/u~�}z�5�<;����f�������3T�ܜ��Qg'�#�u���=��cc3�T����~2���R������t�MbWv�{���gj9�#\�&���t�=+����+��	�+�g�q7P&�g�E�h A�޽���H[�֯�H7߼�Վr����q?��oii�~�j
"bk���E�Y�i�{���0fD���h���
3����H܀1��{��$f&�������*��.V��Y����;�����u�$��/��>`��8D�Hd-_^I�ݾ,�(�4djK�2+������_�$�58A�����ӓO�߹LM�H���|x�{���S*i�����9�X�!�:2�*qi>g� @r;�`4��$�݈~�#�IMTKF0�R�ڔ�
��	�ѧ�1���L�����Z.XL�A�>�&z�[��OLЎ����b�j��}��6n,�|�����}t�/���ٓ�b��c�${A����
�d,H�l���/F�1�N����u����D�YS�\i��"�)�MNy�8̙�o���"v{/)A�����F�D8�l6?�I'O���-B��gt]�jK!���`J\�pXgOGc	���Na�$�8a$X���v�2�|48�a���/��fg��L[$bg��!;`6����ٹ�0^!����l���6�WjI���е�N���؉���۫�~�Z�{�<�b��*��OR���ˉ����+9n)�3�M<�O~�V�j,�s���WR(�N��?��ٻۭV>�UZ��(o��UH�D��m0����L$d����0q0�r#��H��Z�9iI��t&q«���Q�Y'��A����|r*�	�➟�H�Ã����0�^�䐜N���z���P("���3������FFܢ�B{���~v�[W�H�2�����8���?D���QJ7߼���,r~ɷ��L3��t��u�sg��ͬ�B�N�L�K�܇Zli)�#G\��Z!�������B�O��yU�^��\�f���1:z�iVIll�9�NHb���˄���˨��A���۸rY����Օ�E�ƩSS���744'�BQ��0�diRk�X��<k寮0X���B	��1`�T}���^:���&&��94@�y�
�,�>�`�?Kb�7��K��׿>�תEE=�T����)&�M����W��裶6[�H!3�5���$��qPm���X:���hl|���Op�4%0P��6UR]]AF}0N�4u��О����!��9F�����%gLxJ�W������X���\��&���Q	�={z�{p01��A�U�Z�<}z"��+JMtw�kǎ����2��wo�6�HÇ#��i��Ij���Dg�e����2��8C�a�Zzh�9�^V���LQ�PP���͖� Ƣ��zX���n�|so�u�7�T%,���������3�N] �R������Y�����Խ����|(�aH�!����T⾔�ܸ���f�K}S}}��,����T=�8�9�����*	���AVG{�SɌ��r:Y49L^2i^��<d��d3��n���Yi2a��&����T06��fi$���"�j�����ff����U���7�5�UWUГON�O��w�I.�?���K��ﯣÇ�t�=��}��1�AH��:��M㱂,�;y��3a���­|?su�k�42kAZS�j��3����il������&�T�L���?ReE �6�0�b	'��Htڈ�0��V��l|J1n�J�=�b�&L��C�ܳX�&Q�'S�[�^M��E�������������̈Eq��5��ƒ���b��c�t��ַZ�[X���׿�X���m�
v�����}�CzG����
�zze�����ۃ����v6��<�t�����e���le��p<�������f$LV�d�z����y�E�����1D��4"2�mǎ�0}�\(�s$�5͓^�����bu�C�=g��^�p�>6:�e!������oy@BU=��4����A�����Ͳe����j�V
(��]Iwj���F�^jeI���l(-t�%v!���v9u�APN�4w�:;��&����a��E��o������81�|�3��jb�v\���32���Ī�mL�R�.=k��%�'��}|__�ڭ�h
��$���攏����:�{|<���T������C�I���A�Uyys%�'z��㇤0mb�F��JB�� ?k濭�(=�R�3R!!D��a~f�c�&f�_JT�g�D;=ͳGfgU���{�X1T���X�2��0��u�=W*$b�"	Yfx�l���0}�3ؓ�9(|ӛ��G6k�faG��:`"��$����ۙ���QݛRŁ�������b[&:tH�++C�"q�o<�p�������jk��#�D�����C�gp��g���K=��X��s��j2����E��i&�`��c�{6����2����gʒm_�R��a�	HgI��0��4.�%\亪�����zH �e�@m�C̕K.�\�E���� qvm�.= �`�v�q`G+�ŠS�\��#�X�uN31�D�%
&��K� �l
z�ۮa'��C'���l������Y�j��ٴP($ق�~KKKs��=#uZ�?��?����+�?	���nxf�UG��� �ƺ<D�����5Q=�a=�c��DQZzLd��ҋ��.�S��7$��oIIIJ��o�Y�'u�?�1u�5KtMC~��ٙ��ebl����&FF1��h~)�ƽ�\H�!@r������;��Fn.�Zr1��GF��3��k�e��E�� f�P����SW���%A�29Z�h�hll�n�!�ga^x��?d���4H��_.6�)�2��	��z	�O��hv>%����.������>�"	b��-�"^�7p�M����e���q�F>Of��<}<x0�;��
�el�/�T6$�	�c���}��D�޳UY�$������q�����D�f��9��B��U�����=�dC���~�.||>�Y0����;+A0&�cC��S>��6<�uVe�W2L��^	��5�M7527�"�WC�A����mk`��	�j__��544DMMM1���PGGG�W��{vQ�\)�������� H}`U�ۼ�$ ����i_�f Lq�#DxHmmm��؅�{�n!��tv*�P{Xrطo_�~�4߹Ȓ�E���Ů ���`θw2�s�|.�&�o.�K�Qss�؎]�v�·tLOO�|Ζh 8�3��i���J �?�����������A��Ҟ=�	%O��gff5���JN̩̱��pbfffd���]�h D>b�G��1��vuu�/p�yN�H#�2�#���+@*rn`���i�f[8�*3�0P��SLf��Z^�tw��{Xm^��Q=�v���g�P;SW�H�+�l��J+��a����#G��&c��
a���u�pG�v�d+Eߘ7�P:�����9�*o�/��i�u4�L����C�\��j������c�
��:*֬�H=&`.e����a�T�C���3嵂��"S�`��J���1MF.�}��p��E[��z���(��?��nbO��m�uv���,��r9�Rc����o�G�~4ft��!�z�!}j/a*L"��]T%��UPb�X��m|�\�l��VEQ����H���=֓*4Y`��*�S���VDw|�����"�e,�ҹ5L#D>�e4S�5��=�襗T�ړO��WU*33�L�)�������	V�Y|�u�UX�k)���<�-�`/iz�����g�`�TJ�|�)`�Bz�8Ng��	��*�1+َm��D�#4�'g�}4mGQ�!a$��b��Zz2�u39��Ѭ���M����hyC��f��M�s��6��;β7M�פ��U�E6we�� ����͌���`;���]$/q�5��2+�
:�u�WV�n��!/}�~�O���r?8�*/D��^Ȓg�-ѿ�����M�����sυd��+_)���l����|��;誫�BP�=>n��0�z�t�&Z�
̠�B�J~�����t;_=%��#�s�{^`��4!v2*-32��"N�^�ڰ��WL�e?�2�K�ڣD�~2���WT�^l_t͛F�4N�InmEX�=�nVE��5�}5F\#�/˹q�F�����İעb>4����Q�j�����&�4��"�����-�zm�'��EX��Z���Hp⻷�/�;w�����$OT���n��?3��4)�(+��Q�s��������T�0Ss9�)���W��_H��Iո$�����c�[(ZGVK����5 =���4������SDG�F��	��1�}��^yI����7>QS�m����=�����|I��X���R�b�d*�N|�Lt��.F�5�Q���)�@Q(R���nQL-��zp�w�D����TDM8-^��<����l��`��Ε:(���uJ*>]�$�FO�Aq���rzY.�ڍ
?{>Z�/�����!'f�=����ِ���7��J�m��KO�6�ȅ���+���&�&'�Gŕ�t��o�C\��z!��62�Rx��_ULtp�{a��`ⰋL����ٸ��eBh�������b����{t/s�QruT�@���b�AfCe�&	�2HE=���B���9<���L-�D��D�nj�+� ����)�#��^Er�]�)!p���R{&��\$���xYJ�76�.��љ��
�V��쬞8�徉&&�GK��Q9���rJ��t�}u���ng7q����}���j!�XE�����t
x�v�݆m�^z����J-'A<�0V�����M�}��t��-��w�P�d]�K�'/�dZ��$:�/Z����/��|�6�Nc��&�/�UM���&=g,w'�;ϙ���H|�J���P��H8�d�C	����2�;�����#h��|�M��C���T�vTæNl���f���"����`s�2��)�g:;'���e܎����T^^@W_����&��C6�b��������d��ɓ�j�2����]�R�,���g
lA"�iS�`H�|���W����u��0eN��M�۶�s��͓���v�Yζ�/J�^�J\��j�dӦZA�;��&��e��+�h��� �O�`�^>[C�	�A�I���Z.sܸ��c����&��ǲqc�����i��az��V��x8#<�͛���	p�.���?? ���&�7�O#�I����\"��aW���#Mw����A�2�@	��ߏ�֭�d�e�f�_��Z������+˅�8�|v&P�<>�n��-�9;e��Z�ʾ>�hz�/�B@�P�-ֹ�x��UW
����z�� �6�	1�y����I6���@T��rH�&��T�C��r3v�vvN
�R�6t�`���u2ॗ6��LLd�� E8��f�9;f1����J�e��&! �/�@8\x����Ɩic�+��ة��7������B�	� f��v���J�
A���	��S�������ﱱd��2z�l�ǎW�$d/��H��i�z{����5tt����b��gcl�%�@�\�j1;�e__�o0���C��n�n�#��F�ߠk� ��3��±d��g?>����qڠ*�\L3����ő���|�R£�aτ�%{&��?��ș4���Q	��d�G��b�Du-�PP�#V;Q��U�l�e$�5�T�ʩb���&�z�!'K7��K/��믯f/�_x���3���Qp��۰�����Vu���� =��{.s���QvXJ��k���@���P�{l�=���pMM�t�M��vm��\���d��3Ϩ��<-�K�����y��9d��� _�B�d� �"�v�l���'?�g��Ȁ$�n���>���c���8ؓ(�������xF�~��>�FUF��� ��+7�pc�m�e磙�F2�Nup��UN��;�Mu'������/�Ķ�)��&;�2��F�O�w�E��o����{�5�r�%�����/1t!�������"������0]|q	J�?�MI�'.h�h5�����Z����{�-lt}�;Y�Gi˖
Fj��𵵭�m� *����_.p���p�h�d{W��@�а.����p�,�^�'�K�ӟnG��q%KH� �r�ݧ�S�j�N�p���XQ$s�ڨ�kf��UԈ��dﲓߡ^���Nb]RG_��
*-5�����D������RK��wU3�|,��8� WUe�>j�yX-��X^���`Mg�O��p.N�i_{m�P���1�%N�Ga3
�ffƸ�e���FP ���mmk�.�í_�^��Ǉ9��b��O���\KK�T���`5<�+p��u2�.��ޝ��&��8�#��v�u�U3A�R�n�b�hb�V��h ��u\��L�O�Mo�`�P�e,��wZZZ�H�ȑWxNU��'q��W&괠�����2*��boʁ�eN�<2�F^�Y\`e���c���􆚨�IPH�"���:�,��ްm��f��8b����kCC}��8Pi�m��0���Ӣ���R��reAV8ߝ>�)sRيD���V(*}�7h���#Lh�,Y�mmU��gzM[UU�uTTD���c����ԩ4GT�D+��ӡ"��0D�1���p�z)e3��%Q���	��y �Ն���Lp��.�wj�zҜ©���\a��g�S;�tJ?���q�i����N����̋wS]m��aC"�u���/ѱc����F����}�ۼ9!Ҙloo�D�Ǐ{(�����ڪ��1��%]��V**�����+���}�k�.*�u��R]R]��s�w��@m�!�ǜTĞ��c�����԰��*w�^s���sx )6Q㡺��EF�}��9�ʒ:y�'#���j�lz��+��˓Ю]���h��؛�`��K/��eA}g�oV���;'2�A?G"c��	�[<�i�lH\�t����� VTL��~ffB����M�C_p�t�3l �1LN�ɡ�S*���i����7Eq8h�\����T0ѡCs�Jϱ�W�}�$p��211�s�����`1ͨcG�Ίkw�dr�nXU7d�X.�a|��z{�t�]��Njڄ�$j` ��F#*� ���+�|�K+n�9q2>�����t���;{��V0��2'N��s:C�x&m)S����n���V��r���Nu��{�wIw���ﺫ����Vvxt�����F��������wPr���dF/a�#�S'�4�$�$w�����Q��7(��ӓ���۷oJ���W�zu��ţG�8ᘽ���^~y��O��Z|��	�:g��|�k'e��@H�8,=g��)F�*Y�1�SU6���Ƃ��ov�d"�� ����&�����	��Sr �e�����68�4MW�����  F���Q�F    IEND�B`�PK   �f�Y�7}b  ]  /   images/9bbf0d51-8956-46f1-ad90-c6ca9bac44cc.png]��PNG

   IHDR   d   3   ai�   	pHYs  N�  N��"��   tEXtSoftware www.inkscape.org��<  �IDATx��\	��Wq����c�{gfgv��5۬/��)F���("�X�+R!"F�����#Aز�m6���]�w�;;;�s��3����w�����O���.�ݖ�7�]��zU��ޫ�^�]���>D��)wb�d�����p8J�M��x�Q��iH�xڇe�3̣��zI��V��ϝX&��\���U�9��:f��h�P���$X�pbf�!oV�+��
h������i&�j�fJ���Q��0��� �97:�bН%)���#F�w����<�%*�V'��z��fs��Qxg:f	��P
5�����i�Iöi���S�o0y�����)�C�����Q��7�{� 3���p��ӄQ�PG�!�U��;�a:�L��	̡�߻�s2�k�2�	�;�����8�eH�<J�Q�"ux�n�`DC&'��`�0\�`�5ޥ@z�, a_V�i�B�=����e����qd|l������E�{:ZW� ��E��{(Ң{��v!f�?Y�������)wsǌ#��q<?�B�%�*����М��B����ᖫV���qz�O�T���L	���&X��^ӖAS��'φ��u5���˵�^�:nqî$��������ݽ	��fI1�M}o��!�v�8�v ����XN�7���1�<�䲻����%0���ଯ���z�486v�3C3��SC!5��jΡ�)�Gτ�1)o���
�}��Q���Od�b�Nʏo`�)�ߦ�eXm�ؘ�.��ߝ$'��F�%�􌏤t=�����6�`��[	�$t"f@��D�If�ҷ���Й��I������^"WXc,!X%�6M#��(��"b�;+�$ac~�c[rK�J���.��?�u�|h38�X��k�R�f���1ˮ�W�c��^Ni&�X.�*نd�K�,AzYU�λK�D�E�
�'=�$uWI/�F�%�ؕ�`)��� ;Bm���:�t������7#}s���D���Ӥ�]�0���ۚ9ƶ��y��ʙbO�g1a��!�b��o�E��I.K+(�ؠ�P�pV"m�M�M�QOjP��2+o��l�4%@ӯ@_�`3�-�dn�k߇���Ͱj���c��H��drVJr4& �t���	�'�u;������Qlܽd���\T�E��P�D#�9�&"��^�	�6U=a��(ڝ��r�Rdx��!���(�</F4j�%�l�g���G��w��[xn��"�V�n�S���,X��1��V�4p���t�&Bv��P�,a��*	n3� �A�4�{�}���y�m�h�#�����(��wt�&Lj,����,����&��6"�/���4�B�p�:[���#3����Cس�C�?ta
��*Zښ���$��S���mGMM~�h`t|K�q�j/�~�&摜]$�;��gjk��,�p��d����#u����1��Z�;��X+}��� �UD��W��u#��`�ܸ_}C#:;��Leqfp��\�����	~�|���R�>�g%���㖲<�2C4|�8�
�Ģ�R%���l��M�%�]�o��d��	��H��Ko�V�5d`]N���ʩ���P���ġ���IֺX,PZ��2Lw�|����@*�&"9*�P���JR����&L����U�A��ԖN�x�j��`�}�v)U��_P�.]G.WRmҏ9T'���ߔ>G��K�_�Z��TFn�p�o�M��ot|Κ� �t*'F������
�h�Q��ф՚��XM��K�Ee�w��9�7=�$�`0�g���<�BmiV��Ό
���C��C�E ��@3��Bx�0>9O�Ε��Y���qJgrg!�2����2S�o�����ĩ��*��R�X���s?���VI�%$��a���vQ�]�Q�l��W~���tn�qc�[����L$�B���-x�bi���� �����N��l ;щELN/m��%1dc*)���'M-��1��b��084����;�N�q��I�����M��>���<�+�&Hsش��%uLل-�V+GL������XZZ�]w���_����'�p:���[m����xu���ɞ�������Z%�����u��O�63���"�m��������ӆ3���'n;�mm�HҶ�c��<r����|5�UV�|m�k�:9!�M/�gf�h�D[��ر��BKf���dd��%���<v6���r��Ѿ��ؠ�B~L�,���w|�3x��1ڳu��u�p���ٶ��,f
;����Rf��[*����,�y��7�=�N݃sS<��������*�F��jIL_�������S�s�\d���=�C��`�LY��>İ�&sCG�_�닸��G������|wC|��{��lY#������S��u̷��3��1C�]�Cf���&Ƹ���?��]�+9��7<C*��$�.�F2M�By��e��/��LF}��9����s�o?�.4ԇ�9��lr�Y?�啛��ێ��%�%Mՙ._U�,�6�ȯg��c�V|ʕSY�T�������(�JkOkR�07V��夻��V�; Q|�t۠�������(��ne�uy�:K~$�����o�:i	g1�⛿�AW�Mi<p��*a��.F�.�ZBg
z��x�/#\X������W/�POL���tgwCڒ���̹_uy�J3�
.�dc����ئU
۔]�)a'.[�����zJ�y��Sg�w�eqxw�4�//���L�d�t�^S�&u���C�꼁w����l�S�P�:����V���|܃唛�*�Huu��S_bWJ�oL��*��ģ���>�V�8�>O�������n��c��ӆ��9!�}��/h��c�rN��li�E׎f?y�޴�ӋXX\�C,���	��I������D"]�������*��thW� a5ľ�;n^�(#��K87�ώ��:� �O3����������o��_�^o�� �M ��������|��9O�L��_�w|���G߇��>bPZ��q�¤����j2#g���`����� O<����0�����<�����u�a2�����MfO�[ɠ��Z���S�g�3r�~����ŗ.���dp䅳��Ղw�z-j�|ph�iF}�� IG{[�̚���i�v2Y�ֆ09� G��\ՅPЏ=�;��{�M7�G��f^A�sYe�g�o�$����h�S7Y����5!>�|�]b+�6̱Cp�������VM��A�0��3���~�� >����} m��8sn���b��S������8���)L.�֫,���R*�Q��b�:1Ad)N�B�ňo؇G�|ѕU\����)Qao��]�z4�u�"���BLȡ���lC1켨���%��.3g��<Bjk�;���݊���T�V]���ZA�/���Gv�3��n��:ë�'|�$:k�djR�=�����f_�x��uV�RM��5�J;l+N�ˌ��3��y�lۈ���Ɍ`f2sy�����I�5��f����u�)�3���o�&vܵw6�=�p�/z�qg��n�^�sn;��XKj���;*�)֗S�e������Z��՗�Nx�{t�5����U�I�����:�d�{�� �E1�LM��e	6_�s_�.���W�L�h���λ������M*]'՜�����ǃ��O�^��
3!�+��<Fj�g�f�`��p�>��>���y��� ���7ϋ�2���5��͠���o	�xjU�d�����u��� �mwh��O�����+���]�;���j�q�����a"�W�Q�R��g���|a�[l�����L}n!Vv�t���k�z$���i�V$2.��mf��VY��Xd�*_T�\m^�jȞ@�&�~&�����m��28;p�--�����S����h)�yѠ���r�U��y+Icf��qo����=Q�U!�Wބ�ZKl�x���ބ��(b�8��owbp` �@ ���Sr�w���jo%��K5��J���ϊ��nI�
�3rE�kz�c]^��$/��Ey/��y11>�CC��|H�i	~��W���Č�]��юK��_cؐwv��ҒB�z%��.�PЇ��y���������;�W�]C����7�n��KM���'�����;W�0艧^Bm����rs��sϡ��7�r���En.^n��b�K�tPn���U�Ea���M��~�-�ު��iټ����M^�b	�������x\�`Ng+��pb�1�NDԫ�-�e<؁�#���'`��m�\N
��3rH�ʤv�k��H����񤱶��v��&5`Xul�z��Y�`��꟫���G�	&/������tխSG�o����m���6e����>�ۉ��4���G�mү�򂊗Y�)�B��+'Fpwo���W�i<w������߅��Z���3Y�85,������\�wp�.q�O�,b|rA}�v�s��%��oO'��=�L���:����?o��}t�h��؜<.�r�!�n/�i��>,���xF^4��r�Į��]��������s�s��ӄ���j���*F��RG��/Z	���=ޗF�u�^d�"��3gǅ��a|��ߧ�[��b�)�Q���(���y���~^eXXYB��Iĭ�|�`���I:�f��+�����D���-={�/,��cZ2�$lq9A,R{%�J*O3o��f��Nb�I��/�^���ȬH3�V�g
>�OpD���.��0F�%-m��T���r<��Ub�z�-�+���g��$p,�[̀{M�E�2�8'��-l3d�	����)�!7R�]�ɁD|	�ļ ����`bb���sI�K�4�#q!�a�h��[o��))ǁ���U���e5妁�H�F(�L@sx�r["6�Ċ������C,�����KF>���*�y���ޟk�o���22Ɉ�a�R��,]�*r!YD<�}����1��>L�1h,��g��D�dB�1ᮤ� �?GDP�+E��H����Vy���R���6n�yЛE{m\�ۨ�.ڿ$J	��9�連)��@$F] %Ag�eeM"�p���`w��8� �)�j���ql���0v�.��l܏�d������.�f��9ڄ��hJ`;ڄو��&8��S4T���`Rpb��,�֗�ߓ�%I``cZ+�E*M�m��J1ֳ�2�8��͕��fH�̢�;�Z�#����q�1b�	qdP�:�!W�Ys�S��80�S6��r�KĔ�Vua.+$�n�@H����J�S�7�'PD�`�DtuH��ƣ>�R�C��� �0��5��T.�х�!�R�M���c1�<u�nn=�Q(2���fB��pq8𘄧AL��Q|�.��7$<��R��M��� a��z�����k�۩�����o�|����l�WgZ�眛�єV����2¤�-�7KOc�.Y�rT9&�N��s�F�2��2��)<p�N��%?�1$��'�T�	�Wc&�N⡗k�-ZoΉ�o#�/�D@�0�����^��-3��p�R�f8�U�9�{_{�F��)���а�9+���p���b`+���ٰ�&�1��ud��S�"�<�0G,�MJt"���@~��^b����jl��J%C>C�����,TȠN�����D��χ�s(��[+�i�d�T���OPqY0V;cKLF��rr�鱁�2�$��	_y���-��,��c*���\PS����G��̡��0�ϯ΅����Ϗ��ݹ�h@چ�G<��S6��YqK@a�5�(1��ӢT��d���OBE`�G���Ǳ!�ɏ,6r���]f��$�ӎ���3D7s�2���G\k%�(G\sav���}������k�f�6����0�;Ov))1�x@���۰:�J���a�r�yC!϶��b�hk �dG���Nd֢ޑ�X*���^�.kE�c��ޱ�d|�g�D�c)ZQ�8��4{,�������L�����a#8�}�t�?��q�d�    IEND�B`�PK   lg�Y�{�" %# /   images/b7ab4f1c-086a-49aa-bc93-bd307c85ad93.pngԻgTS]�6AEzSi"ҫ� ҤK	�H�B(n(J�4Az��PBQ��	��PBM�oo���w�ߏ��0` Y{�=�\s]�֚��}�K9/B �KڏA ��j��<�I>w����#?d, �9c�Ø|��n����u�J�z��9��8Jx�:��)sB � ������M�M'�RYU�xb�$��U���l��KƘ�e�;$7S'K�&�:�������y���j�P}�������S@�z�$t�M�_~㗸v�1��t�����4m��5�e{�j���_*��_v�D0���ٯeQ�0��%���>��K"�K����PAn$�� �(A~�dI�E|Q�����E=?��C�L�tF���!҅3<��Ǐ\����]afn8
��JS=9�~���ɜU�Ν;sᢼ_���SGa��t����>�ke�����oOoq*��8B ��g���[L��_���vD&�EED���	���z���S逧B��kj���ʺ�{��Ęl_V���6�9��숞���	�79U���-ok���Ϩ�wR���2B"|��i ߯��iI uT3�j�d0�QpŤ�x{�Y��U�ɶY���#���h���Frǳ����$�!gr΁Ơ������}�k����}z7���D|Cm� �.��W__��<��΅��߿5GFF8�����~�Ka�!���No;Ku&)9�h�y�艓S>8��.�����>�+���$,��f��Ǖb
��ϦYZ�L�����R�TD%ʇj<GDo�~j��ƄB�3���ם9�� D���"��M�>a~M���g����w�dƆ''���*��m~��9Qk^RW�o#�Qq�M�*���kg��e�O5�8gN����[b̽b?�q
Z�6UR;�+��534$��v	B�r�Cw:q���������26�������(���ʧ��ku����t�F?p(t���u����-�vES��S�UOc^YK)~�M��d����)a���d���d���t�
��
9x����3�Z��a��O���8LICex�}��j�I-..>_T<� �&��yu��ë{������>��it�׬�/�!�o���TN�g}hO+�D@�Y��8�H?���U0��b�˯����u3y�'3�+Y���M�>I).��|a�:ϟ�3�L��В�������2��-����e
gQG	�?s�Z�k�>���W-��7�S�4����Q-��zep������t��{;�flaAVe�3�<�X��j`���^�J*����d/Ҧ��8�؇�VH��>��T�wl��;�{���?f���Gd_I�[��h�ɸjj��¾�~*o
x��O��n��ݹ�ۆ��f�8 x�v{��!1�u�%��<��7呹>�fED%����/\�N�Լ�b[����"�b��
"u�ƹy�v#}�o��e4��P���0L(�]�`�_����W��~`jb$
��4N��
\v����c��%����[[8��w����iG�'��UTl����(S�,W��CAX����;�CT���r�AE9���uY_�<�вi?>��_4-!�.hƨ��-�\G�&rH�o��pAfy�<��.����n2+�i�.�e���������~���R~`F�ҙ�[�SR��l�tAC�=>U
��	9l.��I���1�\����8-��V~(d��ѡ��q�$,�;�Tf8�_ �#��Q�NS'Y�6&��t��<j��V-hIV�SO�h����N
���"�VM�6�|�uӐ��#��(����4�w���77L~��8uvO�C�BZWv�'"�����)�c���#�ۋ��D\I��p��-�����-���b�x�B3v�*!;.}_Tp-�-�++�	F��U6��CT��&xX�3#�����-�dҽ#�YVܪ�v�`�.r]������uQ����_Ia���zRRRqyyr���{�Hqz:w^��s�$
x��!z�DF�$N%�M8�h�/�-��u��b�����>�)*#�K0�/*)i�ji6i{+�	���n�*��aaaQy맽܄kD=~��E�&�tȎ����C)�^%�E]�&x��+��0Gguvh��`E��c�E��+o�$�@�U������Դ��>��::��D!�0�/�EHX���9Lq)�r0i�֎.��`>f�c�3iѽ��I����;a,�VRH�!��K����G�ؒ�� ZQ*�}�^��_���Cȏ���\ء}����7�/��B ����n܉��R_�K]�E���O��"�c����h�l�
*.|���EK�rL�!ny�7�=�t�O �-[�GB�&�@<���(qh�x��r[SC�-�w|-]����ݻ
�9:¥ȶ�a���A���7eFʁ��d���XO�_A*�.��O�[�B����0��U|&��_t]�1��)Sv7���CM�}�o����''>�R3�����s�d���z~��,��ȶ[C�ݺ���3��	C�ƾ��u}K�@��T.W���uw�j�OK��aL-����/ҥ����WJ�q���׏�j9Z�D^�����j��<�"�33�9j99H��8�P淋\\�D�)��O#�;z	�U�M��~�8�
=�z�<[���l��H�((-����9��b�o���'&��_�=K�bCL@,�CK�G[���F��9�

�&�����Ώ��e�Mߒ�\�x�Pϔ��8������4���=F����Y�F��K�A�Nȵ�Xs����8u?�lG+Bm��8�w�5���~���p ���Nk����D�-r���0#��]O޷!�F���C���
�E"���$�K���Fn*�})����9H����w�,�w���~N���. l���iI�>���!���M�|h�~@ih�g�)�f�� ?w7�Wnú����wܳ���G��/�L���$~�^��y�濐2�A��F��D�J`K��H*��ϟ fu�����������l��D��L����ͽ�������W��G�gc42�,˄b�9
>��V�����饽oi�tL�AVn�i^ާ	\��C�/|2��u�Ih�Z�3����Oi!�7����%g��ځ<$�����e}���� �p��+k&���[[=���#r�����7���<�ݍ�o�<�2��23%_���_T]W��H���--&%��OMO��~�� BS���ٿG�})Vi����CO�L C�3UZR�آ�S;��\\�� ��k_qSLD�#E5aaa��L"������<�3�����7��RR� :�����+�����s"�ݙM����߳c��o��w=95d�g�2KZNM�_��>�\��� Yo���R�'�q����&o QFذ�z|V)�1'�S;���?�N35%�7ӯI���*n�BUw`�ǴĒ)F,Tn�p�F�O�P��g*�?�Zj���żi�����&!q�"�pizv'%13s� �mll,c�3�z���_�Π�W��C_�tIH�0vp�-��j�g���LR�>@�Ѷ�.9]Q�N������VA��j�EE��2�.�x�O���sBz9�62V�`
��uv>��RW�{tvtZZZF�������O���ĩ��IJH�'}�T�`�&o�2<������#��p�``OgW�	A��;YC�o��gQ���J����4
ƀ~��Ο�!�֓?7�LPH���]��]�7n����r~~DT��:M�v���LR��Y�Μ����ub�Qef��>C��Ә���ȹ��Ϩ\o�76�q�s\&n�`VlT���D|��x�������G�edb	dIW���v����Iii%��f9:�����e��\C�4�'9�
$�qE��e<P�3hD�W-; s��������t�ɬ�s[D5̶��߿B����O=j�O���\���_(�����O���R����>�k�J�4ھ�a_�U�\������O�hk��C�1�),�#б��b^~s`$0��;ak�f�{� `�Icp��Yd�v������Y� ���Fb@åR�k�����
~�n=�P�4�eKd�E���DOIU�?l���-b�.��Q��Ț�����peK++t�I���3`�/�Q��'o>� �,-δ�ҥ!? �D���L�!оtI�͓'�1���,�Ⴆ�
{��O./=�q��]����E���Ş�cu��⁋�9�LǪ��k����33���� :��c��p���6#Oܺo���-%^�-!�%�P$׭s�84�LWY���X/:Ui���s�^P̻��w�r�6|�E?<ym�ɟI��o[� �����==�_9�� #ȩ�1��<<�#i�h� }J9��E���Vl9UGN�P�ú�Ф����%zڍ��fX�ϯ+�gT�[�9]sd���Λ�j���O��J�5d�_�}�G������`((�	�N��Vǿ�u������Z��w�] 9/��3t�f��∩1&�c�xwz�o�w�w�89�O�*#���uُ>����+6�@N�<���t1U����I���9:`�V�1��iF���6��������Ja^_gs<s4Ũ_���pr�����޳�D�\Qy�#�CC��j�7�fn�5�ɲ��
�H��\)Nx%l���T=��k��c�Pp��(�7od�Qq��z���(F���"!�4j�#q]�qϩb@��r�"HV�ITR�7gTd��k������rȣ�(ʔ@>Fa"�w&8"U�YXzpt'���j�a�#��S89�
Շϑ��k�B��7�M���K\v�6M�ԅ�� ��ds]��}�e*���>A���}𱯮3}�Y��{
@P��
fr�T�9��̚L���L>>��j��h�h�gA�&��;�u���8�{����-�r�n��#~���Yf�����R��<W�(H �==���'��F� Ci�3���E@8��	 �E��|�js	0��1z�Q!���v���J�� ��kG��@���EHh���� KO*�9«ɿ�L ��(c��(4a��6r���F[��.�x0�@_�2��������.��4��p�D15F���%ٵ�0X���A"�嚺n5A��PV="������T�t)[5k�Q�S�;?p1r�y��	ЋQ�}�U%[��&4�9{aa�ZVixާ���������c*Hv��-�[�!�f�W �ց��S��lR��O��P2��'�e�K��ڠj�{��^0ߕil�6M0�@�M�v�L��=u�cdUȉ!E�"^]�s'M�%{5��9:�dd�,+f��t�6��
�/��Xڹ�Ga��Xr�����g���u�M��5�~�2�vᗮ:27�$����G+��s[���e�q�y��6���s�@�u&�3x���Lt���i�@���5f�3\���8/vn�P�\��0�sbv`:� kDԏ����ڢ��#�*��5�{�KK��Ԋq�1+c&0p��Pb�V7N���-wI�����u�nD�iT=5�a��۽!��=�����gj�r� �'��-�ֿ5_�U!Q��wIq���EyU@��&`�K���766_��sm{�{���(->|n����%�>bu����mL�+Ug�n�����~&�N!�H�hUx�穄Vbmx��ñ��Z���a�B%v��wK���Mh�hV���N��+#nS��.
 �����~Yde{�|��懃�lKp5�B!�ǅV̇�������vv1���<� �֗�9k��W�a���x���=P��gI��lX��tx��;�d$v�#ג�:��G��� v�O���Y��]��w��P��Gj[�^��/�}����2�� �G���	���w0�a�����Tsx��y ��g%0���E%I��FPw�P�jҘ�(u����#2a�0�&'��f(��=�̰8�C��<��@��A0��ɯ�%�u��q�Ȱ�Ys�^j\sFǿ��S�dO����^�P�V�6�Jb���	�z�0�=H�����o�/���;��'����t����j��+B���}e��%hU�iԳ�
z�������,Xzxa�<R_��*4�1������*�M_鵁�Ԡ��>`!f�v&*��������E]]o�eS�%.�-E�)�Y߶�����5�ⳅ3'K[����`�R Ӳ�rB�+y�6S�,,+�es3��Y�)����9�X:Ԍ��~좡��c�*2T��w�' a�0��ҋf���#ϸli�#mu)��F���ݾ*�NTa韁��C�3$@掰��a�e�F���RUޛ��e"��6PZ�|�F���/�O �0{*��ZV�|`���Y�r���������KP�iެ+9q;W:O7�
kF�B��L(��E��3�N���_q˻� A�t#����xe,|���j]��gLw�j����$���x���ҁc�'�j'ܑ�m������c	��^���|�87w+ ����q�G��Y@R�*��?�D�q��5`lBڕ�j�P�����c�����*���%��"�t��%X�et���9����2�P�3m��*5V�M�k�QW��S�U����]�W��B��6��b�PS�@�J�y3k<���M5�/s�eQG��f�J�o�O(�U$vv�����!��Q�os�n$�48�s����5R|��
�V���jR2P�?~�&%V�Q��^4����;N\c�*�\3����3����?���* �B�tv�ݱT���&W Z�@x��]+��@=d��[�
�L�G��ۼ*ܜ���ᄞ�@��i"��֧�4u���IV��� �������HX�X��zyކD]�/P����Fq����XOT���G��I���翨X��u,�(���B+�	��e޽#�"����V0c���͛>vy3���6(��z\���e��ߟl�F=�r��k���O�'�g��߽�%���¢�Kg�0�?N�gQ1Y������Mc~����1���qO��5�}BNi����<d�]İ{���W55EpL:�Z%��y�������39�Ù�f���#-0,��0��{`QM �"�e/T�Ut�8=$���2�+���Ph��Մr�C�*�V�2o�]{�#��%��`-�+� �c0U��z����Z���[/�NV>oS___���v�������z�}��ۼ������� �����Ju�@E�}ɂܞ��|a��G��9M����������������k�g���|2�g�3W�,Sa/^��m�k"!���]��EEevm[2�SKť�����.F���TmD�7����n\��S�g޷����k&��כk��=E�J� ��K!�[;kk3
λ��Yk��ShL
E��-��&6͵2#g����!��j��� �|뭁o7OOSwww���{Ѳ�����_����ǜ®͍6-;D�'��y5^e�r����L�S�:�a�n�e���6�2���Q55S�d������yv������ё�������.�����{��h|�G�e�D˂������ң��d;���ů�B"**�KKڜ�B��s�}Sӑܦ1S��:tx�r]����X�ֽ� ��m�U��ܘ&�"t�,0�eč�&������ e�k���˾�׮Yܢ����u�X�7;�����ݩ�!}�u���I���A�t�{��1;keO4���������_[����q����P�''l�WZ�\$X#)^͋�u�J6BW?�@Be���Hgp�I�mnF��1�3.Rtlnr�9޻�|�b%io���ʉMM���]�k��v����!/>~G+r7(ak��憝���x������1kUO�6<����gfU*-U|���ld�~����p�] �r-��Z�����2��6;%��WO6�����f5i�9��d�a�TT�-�]�ZZ	Z?��]ͮ�voQ�������������`�c<�k �n��h۠0�Գ��_!�������X;j�O�[(A[6�P_�P~�ܛjjh��mYo8��O��?���h��3�W�yj�P�u���답���	=�*�r�DH
�qs�����V��x���U>e`����O  R�ѱ���SǄ��K
jky�=jvʏ3Ɖ�u�j������[
a�� V����&c�͍�����33�k��3߯���(����Z�X(ȓ!ߟ���=���+�Uaͯ�B�~> 2�b6X�`�*�V���O����@��V<o�i�U���vy��=��[���E���%�Seܓ%7��t��E=���@�?����ݜM�򥼦F6)1�����K�ܹs�2n��X xm�i{:�[��Ιe<J���~��bfx�W�T�	��7����.F4 �c�v�l��#L������RtEo����,�I&DK6Z���������/ ��^�a�u�����x��'$ ԕ[/S��z���q=p����@3b���;46V��	�C5�XF�P��4�~����x�dvj*�VQ�l�"���֓�����PU�[�9]`��s@τ������]&��9�_��6�щ�����kaaa�?��T�	X�\�ԓ>m�.���|z��GO����J����Ƙ������m�����,����g���St�q���z�����|g��	tx�v-��V*��>Jbw�?�4�U}}3}�ط���-�������c�WY�1�M�ڟ���1���_WW=x�7��倀�;w������1���R3��`X���:)�������Ń�|��lIe�ݽ!5(����Ȣ�u�u$���tI_
��e�&]{�zr���w��a?K9������ �k
����� qY�[ *�;6*�+�{�L�H�	�`�����eU�����흋ۀ��tޜ�?����Q����������_��"���4)ɑ/ޝ���s����>iy��F>�G�Z�eg͟�׸9�|��U����XOo�5x��Kg�����Y�#�p�6��h4������͞�%n������Y>o�k�v����=���/A�-�!���/���[`���\�%`��**)�6#��r�x����]iic'?
�^(A�'��my��&o�������_��=���f��K�\ Y���*#!��W١~�IJ"���<ZF��G�`�m�/����+*�n���P��ֻ�4VSSs������_\�_'W���=�Q����qG)C��+H\:����1���^�E��kY��-�T!Ax��������9!;��2ZxZ^��B�/h"/ -I))"ѿnh���3��No5=��ڏ!2��@qxD��p�Z;�o���ۢ�I��\jGH�
�`�t�'~��3���5\	����Q�66�}sss�:�|zJ���X�������###��4����t*.R-�Т� ���;��i%և@�ײ������������)�b/��-.-]x!�Z�r�����n�������=}��[��Śq_ʁugj�RRZj���s�<J#�� \R����R�h9���bZ�4�t�������Ay����E��=�##�&����: �*�����f�f�]�+g�Se�B�dU�\�?U�GZǡnn�FƑ+c�:�y�� =1�]��� ظ�WVU���E.w-n>2�ו�\�@��H�V(�fQ�v��	0����щ
j\O�j_�ê����9��K晃,1 nf��m*^p����ԊJ�{'<���=��0�<s��q���j�7�%�d��t<�cralJ�������G�ID筨��E欬W�{��g5w<��e���J�{-U��H�~���+�E�RE
X����z�B�hm�PY��9��`�߭k����7N2�BlSr��7ͼ������}Q���!Xȏ��e�a�ܧ@��>�x��p�J��첺w"�������F8H�g1���û�_7w���Ɍ,|�u�0�=�����9�"��[[[�]Wo��4lmo���4Z�B� 	e�N���v������u�����o

�h�%�a�������:��%���]y�hQ�!H�-�Γ�.���ϟ�/*!@�r�kG� �\__��ۛ��ؓš�ib1~<VW����N`����	�"Xu(�~|(!o ��gw��ʕ��[<|�r��� ˳s�e�/AAK�����)��^�_�T���'�������i�fL<�?����F�(�'AT�C�h���+@|vq{�`����"��������D�����jN#ML��/��TLN�|iiITD�PC�Հ�u�ϺB@~QR:���>���2G��<7������dbU��GE�� ����
���)�+|$F�q�I#���"���wL��@��~��v��? �q������	$��P�kL�t�Y�J�Y����V	�ڗ��L1&�-ք���|]!c�Q�J�^RR���p.nyW�ji�2�Y%�	%T{�ӏY��>L0CMMp��r�c��Q���j׿��̖)�*#���w]��++�$��d�ɗ��M� ݁{tU}^����n�Z+��3|��\g��������J�FqhAľ���mf�g��Y_`ż<�{�L��흗�{);:v�� Г��%�]i�����!�	3|�
`nO���p��㡂�P=��᪽a9��.�/!^i��+�=��c)m9�v�ׯ�)��}�G�@���9�iaﳊ���ט��K|3�!rF�&�ȕ+{��1.5Q#2�zS��6��oGU��(��rQ>��y���K�n]Rځ0������r8�|4}"?|,�;��|@�7)v&�*���(p�_��/#�C$y&������+�c�����.��v�-���#�|V
�5+è;���	�YO"t������"��{�������2b��l����2$�蟑!Sը�>��Q^��F~X�����8��С:t�>#pJ@P�����G��ԃYØ��i�:�ڰ��m1���껑�C<��Ё�c��>�l�Uc��_��E%�Fʡ�n.�G����'�H��C�0��v > �Q�`��}Vf�.�b��ъ'�@Y��
���[�*K\�9�d�4�OU��7p�|�/�8��=�'m��GB۩Ji�h��3XTP>�C�;�l0���=o�z�~-뷦���M��\�R���B�q7��Kra�x�xw�Zxr���y��$UA�����N�N�������E͘�3�Ҭ0���~P�;��\ڶ��|D@IAl��%������_�����_�g��u6���z�?ݲ�J���`�	�=ˎ�7#N�EQr�����E�?�R@��p�0C������Y�^�s��uT��b�D�`	��xA�y�Ĵoi�����o.ݟM 5���h�:��t��L�}��_x!#�ý<�;��h3j�Ԭ��.>>��բ�1D��k��8h�6�1���	�L�_Tkɛ�m0�5����x�n�*.&�F��<�O��l�
���*���g�V��.��`���<�ޙ���F�������B���C��=��+x�ִ��x>��;�y�8�h׎�US5gT*���K����W�4A�����lC�^��~���c�>	����kk�o�?9��������4X��дU�;9�ߑ��U�_y;'z���w_�f�ӯmQ�
��Qܫ�4�S��YA��n�l>֯YyI�uC,����Y�`G����ICV/˖
��QC���(y��?}��j��1��#���R�Ъ��������
>s'�T <�aa%���8�����0+�*ǻo���q���ͫ*�.}(�zX��� D��p�aV��򘢍�P���1����M�_#`�\}F�RS4����i_	n
��M^�;
+���c�����J��un����v�~L�u/�yW}�r
����:;�����{�Vө�J��X�u�`�<��ߝm�|��$�U��5�Hs	�������a[	�%���i3$+��/�
f��a��<s=�:eZM��ҫ��Ӳ�R�H�;��2����[sW������צݵ���WY�X8#�	��>2�)�5.d�����+f{!����B/�HQy�-�m,L.E�hY�$R�tD83�j�;�"\I�侎����,�����q�&��m�a͘�
-�;)O˚^%Ե��.X�`z�Π�RC��ɞ��_����XSx&�UF5��?�o4��~����8G3�l-���?N�����9e�2ټ�����z�l9m:�x�g�BG'M��dA��	=���H�D����N�J/];;Z.~�m�9:M15���v����<��K	��/�[2C��8ZY�U�J~�H���7^�t'�`��c�쾷��R:>�j�Im������Dfԯg���t����`$��%�8���1 `�v���6�� ��������F ��BJ����)6�FQ���,p�^��ɶ���Q�ֽ+�;;[� T��;δTC��֙fa�Q�ar���e��v��m�������+���$��W{���X���a�vx��'�)�4�`����u��yEi��[.�،��^�`��Xu�a�����f]��a<	��F+�ƶ��Ľ�I?�Xҿ:z1C�/h�{�j���t���
Vvɹ�3��2�E� �Y6|�&���!�H��\�o��E�Ӧ��>|	Θ
kx�0�1���#�oU�sx����!cNа���D|]f�LW��b�s, [}7,�з0:x���*�o���wg�����hzM}+��Bm�塁exB�i�����:h��� �񊋎�r�L�k%��uB����$���!��I��J�����<j�ήש=j-V�޶�i�c{�)�5N���C�<Z��)*^�(=�S������S�Q@@�����r��3K\����ѥ�������'^�LF<	8��Ч���)�TU����+�����Л��{�a�O IE^�/�B:�VF^1�)�[|xx��Q\�5P�:`\A^�鱞6��()�kN��WZi��w��1Kc�_�xZ���[�WZg���?�{\�z�� �0����,��(^Ƞ�3�R_a�1��5O��b���'@b;׽��x}��hw�!�CS��FO���O�$���c<Y�/}���ra��C��5����$����F!t�yH�	��xe��9�E,v����<��]�RH+8�s�[�
�Z����b��ǰ�-=�q���l{Aคx��������V������%~<�-0���P���!G�H��,qpgIcv�+�� ��M����m����*&H t�O$�)~@�U��uu��E�U;~�;����k��u�.֘�OZ�py�Lc�yDE1��7%OR��aKU}�9����F/^$$K!�7"� ��)�@k�]�#����q}��$��W���WTHc-k���;�-�ӭQ������(� !��=R"���';X!쌄��˯�h�u,��.��'N6�$1���zS�h�2O�귶إK��Y  K(bjj�I-���KP�ZZ����-:V�П�>A���+>��J��:y�Y����d�`�x����Ie����x�+�F�ªjH��:�}:v%i���m!���5��hw֯�l�FCm��j���L�+�:��&��0��5� �F��f��79��P��[W�m�]!�����������Sjl�[���vR&��I#'�~Rq�J�A�L�2���67�c�j&�3=8x�%��_;Q������h�d�����q_����g�2���!Ҙ<�xٚ��%�'=%gihB��η�r���Ke���>��)h�3���������]�b����_Ԥ������OU$�K$�B3t��zZ=���ܮ�XT��w��U>յ��	��P�-Ȩ��f���Q���W#̠��բ^��o����"%r��e��i_��|���e� ^�L��K����%G	
��%�-&L�����o�c=�],���qZ���h��+d��fB�Q}Zy�����ڂ��'d�4O�趆p�J��,Qq�Y�:�;���F�ii�-� x)Sb`щ 7���'<���K�)GtKo�+�;� ӳ�S;�۩R�o��O�x6����X�vfK�؋��k|lΦ�
����c#��e��'S��nnҸ�� .^����3��*�@*�V��&B���¯�)�JJ"����K�%̑Z��mK�����>R��OF�u�K��Wr 6�.Wv�4��X���w��v�#�,���R�������.g@NM��� 9�ܼ��M�̱+�����O�r�R�rQO0y�Gs���]-,+E��%
Oi	yL	�V����23)	 v96jbb_����ڡu��s��8�{ߛ.	���\��'�۽!ٰ���\HI��V̗��9]ۈ��j���� f��Bl]�_�!7���C�vg�� }���䆖J�Ҡ��b�+��i���K��O�l�>�o�	%h� ���f����4Q�ϓ~>Hs��-Rњowo�#�;%�'�O�U���٨<-E��Noá`���p�͑5��N��؟��E��q�l����1�.��`��)mn��p=��e�x��)#��������E��8T�}~^peg�1����R��EaQ�]�t5���IW�U�j����w}�گ����RM����o����˵��>++T�/���͞��o�aZ���4C��x�ȜV�3g _��A����r��MTN�̡2N~�Դ	��)������8�,�����/����>��<T��H`ˁ=���K��}��}PY-��bT�d�[��%�0��L��\ g��؄L5��a�與�\r�]�����D�C���}�����jC����I�!�sH� 9��n�M�5����׊�S�)U/�ʖOp�B�XG ���Cʱ�}JF�-��ܝo� �l�s�m����:g�H���GO �b��� �:r֔����*��}_T��.�y)����uK�w-��+���	3�BC�˞��x�������C�ӇR� ɒ�Q �l���V�=?���-�F�M��!X5�%�S��Հ*e^!��f%�a��1��O_�? zO�y�z��7Ň��[_pJ� ��kUw�L~��7�0X�o-@��-�j�D�jhP���W+�:�825�@���M��X�B�-'G��akƞ*�݀2�g�bHK�x��P��lL�Y��|����%���9a]���@i�N��W�A=����� O�� ��6^��<>Z�12L�6P�,=&�t^J���0+36@<05����m���󽱙��bw�-R8�S����j�73��������[���22R���>W��=����5�9\NR�t��*�_E�t9g
涥ľ�`��G%%�Vû��K��|����gc�������r���᛿�I�|-�cv�'r��8?쎆'�����
>D�=Hi���4��9 %2��@���U�^��(Hh���NQhE��e�p�����j��sQ�7�/`0��$������|[BP}�m�o��X.����C�ڔ��؅��G##��+of�j>6ڳ@/ޔ �:-w��U>�<��^Ό��Ǧ&����.@������Y��ghi�U����r[6��D�9w�#�n��[���1:0D*�"ֹ1Z�8�k��_xW�MVh�Hv�M_�,�U��<J��mx�LW�����o|�@5�髑7�ߗ�D���IT�V�J�m��
h�_)�!�9�m���}���rb�>�{�����;iz����w�����y��7�''�O��Ց$c��!���9�I�ϰ?�q����ؠw����[�8J���-F�.�{��&:����z�~Iǋ�S��}'�뽳������^�*���4A��������_�. 0�����	c�m͚c~�����4�Q�c̱T�:q�~*�s�o>�W0�?O���Հ^�X�^��W�Z��}rZ��
S����P���nl��b�l�2�ķ�}e���Z�R~�{D�A[y�Mf�L��4����񕾰-�sG�0���Jފ��t�n[�6!G-֕�:�|@9�j��L/�֗�N�]�2S�hxAiX?�<	e�a��'\c��(�>�stodd���<�c4S9��fy�1�%�dt��gwi4��R���
�?!SU��q�)k�p�Q�WKq?r�� 8�lQ�<4[��dۇ��4����l'���h,-�μab���3�%�̊��J,�;�䒠����'�yT�m;�+T;ٖ�;G��U<��4â�w�J���! (����ố��|/B;�4�B���!�E����m>�;?_13�����I���X����0,����d���	�:�h��Q�7�qc��ּ�
Q���J�FǞ��84�w�Oh������4SH2�$RM�]�hp��S�7ay�kzl��|�Խn�@�
S��ìo<�7_(|���[�ߎ���vm�܇��`�*i\�6�E�h�v�j��L�M7�u����I6�a�_�wf����F���SϺ20@0��׈�om�8�P(FH��
jq��Hp��d��ӌX|q�����Ғ:5%�z���W�6Ѳ,A0P}�<��Z2l3c?�Y��sՍ���	a��jUG���-Ɠ� K�b�pF�޶�t������ͨ�6���p���Y]/L�W��~ޛۤd���g����|�/��]��������a�S���'yȞ4󖓱1�����?�B�֢�A�}B6N���<�0��W�1f�x8����j�����~��D�W���K��,e���L����n�lll=�OmZZ��ޕ�q�g�=�B�{>��?U�є9�v���s�������=��/_:d�Y����I�-D���;b2d�ի���F��(�N�n��ǭ�����Z55��Mm����2,��{&�%$tD���AAJ���F@������k��������>�ߋ��s��י��Z{�{��>���L�K�WdFFF�IL�Ϸ5�]�7�ۿh���p	S�wS\i�W-:��i���w�\Fj���D�����������ov����,��C5�?T�u����V�j�lW���1������^8�iR�'2t��y�W�:4�C��?t���y~Ǔ7��޸� (�dNW,5q'��=4��SS#Bg:�Uį�,HK��2��x<�G[p�����He���o�4�\�l�ނ̮h9k��=�I���W�[pu���3"��,���ZBaj�^FSp�R]�<�����<�V�CZ+B���SP]n���]����7�[����0$I�]+�KF]_��*xt��ˍ��J �q���$�p����M�|�����=N�t�,�(�Y�R�R1�/6����?5u��+�J��q5lW{�{��~�p�ƹH�%�Y �;��/�c�"��H?)��{ha\fy����yDJJʐԧN�z�SRU������U�ܽI*Fi�;j���a���o�<C4��ǓW��F+e���[�
�V,%�Hy�h�uu�洋*W0}X��WU�WWW��+2&��*�}�������<��������n�ї��m��|8����V^��L�]sO��J����x�5gy=������y�_�2IN)W\Q��𬱧�'BdTMe�l��a�����A
=��q���%������D�p�uK�~�c�.�?�9��}����P��]~�P �"�wv|�Ɛ5ջ���P���ͺ_��qg}x@��ڨ,�{�y���
��J��w�tX�.�[�|x>�z����$\���]�����&�>�I�66,DvF(����.D��d6�K��� &4JZ<�]�j��5M&��	Y)g]CQ�~��%ڟi�^��B�K3�f��9�����O2A{��Uyw��]���駩��>$@�ν;;̌�H�k��$�����4��G����9���N:%��[�f��']݁�53�a]]ݲȕ�������zD�vlҏk�8�uH�{p��J����_�W�8(2.����E�c��l|t4�y���?7�������4���;�)���Ni�"V؞���vR�ފ�@�Ü��+ϋ/��2h��/WV�9	�,�6�_������I�#/�lmTTĚq��R���*E�P%h|�A�\<7����O<w@��ғm�(i<����N�,ԙ'#�[�ߩ�j��O�����Q�!��2Ta�\$���abҧ�	�/�8����Qҧ�ꊖ{��Z�����> ����?�}����r�h^&�/�$��KJ>��Jq{�/Z��n3g~rb���^p�wp�7�����C��V�d��_Tũ����Oˍw�t퓫GH�{�2�@��i �IN��k|8�)����{�K;;]Xs�Ӑ���zu��wo�Ǫ����!S���T;&����OZ/�PA*C5����#`��Q~�u����-�m��}��pKU���Yuo/ �Ko��spu5���݌
Ċ[ ���-=d��UBa�Y���|EG��C��^t"{OG� �ZR.��[�oS���q�|�G��0>#�_ѡ.�y��c��a��&J�����n{l�ޛ��:�����P]Xh�_?�v
�H��*��xk�m1󿦤�'��}�1}��L�V{������/�8Q�>g?3�E��}�Jk�Y}��ղ�+n�1����xP����_�����1�Ѵ뇉�D��]?)W�{���}�?�Hʣ�J'?���efa�=�R�$�;WP�27YaCC���NKK5���y�l�A%�����������ΉH�����7e
�0q6����A�ᱛ���Ӣ�&�����aPcjjjJJJ��RRg��|��>��|�/@ �.n��0�l����qW��������ҍ�}A9}f�W7u���V}�T��4�& H������0����pGoj}�!׾.�X,,x������&{�4XQW7��e ]XX��������T"��O�����ˊ�XB���jaa4^4���A��=ps�L������*�7��c#�=��]=>9��S�.� P֥�PG!� T�1��k6���W�x^�5�g4��8��̭�p_Q:K++���n�-�/Q%Q:&��Ǒ�L$8��$8��?sf�x�*�MMMz��ҿ�Sh_.�wY*.�0Q'�+ ��~�*��y�����CaBn��z>��A�B�ڬ�-5�}<s�	L���8����4rqI��v�$�L̵���؍(1��6�n�H�2�w��q)[��b.�M����~?����6]r�����%�K�s�cy*��_��Sl��4J\��*(Y����V�[LUfdM���}��]צ5����jv5���l��iKKu����z���c��}}�K��Cq��	6��ްi<]/TA��q��@/*j���1�9z�T�_t�ϙ?���i�w��e�����\�'��c^��C����ʃ{����Q �����Vf:��ޓ� �=[R8�1��,S�,�lʇB�VG�t������w;�[���7&ќ��p& ��A����X�Ƌ�L**�|$5�!yB}Ӊ'dA'M���G)�C�Ź�u7]|4*�_�Y��=�w�#F��4�	��J�(�aw���2=�1�Ɲ/u��-��.����R}y��P*w�r�a,0��Ñ��^X#c�����m����ˬ��Wgj��R��H��Eu�g �qF��������ꓯ����`Wj�㔞|�t�~a�,!Tz��γ��vln���ƝgV����>rH��B�h�G5��lGO�F�ϽH3��M�s�p7UT��ChE��.~�]/��҉b���p״-��\n+�B�4�~=YA^_A����t��ƺ�Ԭ:�%#��*;iDL^ݕ�v?=C�5����$[�l9�*K]��������0��Hk�����?���_b�@`��?1nt#��@M�ս�3%9	���E�k�3TZ���ɳOȇ���U���m���Ac~�Z��w�^�@��)�[�����hIН?��~	���Q��}>��p)�z�"R]H�3"zt�\T\\RR��Lv��Q�@.�JU<�!�c�]�V^����宯t�J��=��o,A���9&,�+����Ls#8-tAGG�1#px�����R�f�}�� I<�u����+�Wu	b���ľi U�/.�z�4~��6��A.%X�'
�y�,i�6fϡ��������=T��'�9T���H��3����PY#6��S/�?�1�q�������ȳi|����ë��8�����U��c��t�-��9����ÈU��%��AKqhg��y�����ɢ�t������A�3���K���AD���I��k'��Q����R����e�<
�\��?)ń���5&����m	yAIK��;����S�+֨�s�i@�G�YS>u��ׇ�Y��Z2�M�Y�!-�1&glL��8G��jU����S5�
x���^��k�����B�$���/���w��P�L�''��ȗ�����✕�T�f��Tx�u�NI%���� ��7mTk��ܯQ�VL�"��"�����O��S�J5#BO%��~C��ɹc��
�BR)��`2�a����h��"_L�Y�^�5>��=��5;�����t��ET�͹��\�xT�ܛ� ��u:�h^/���]K�&��,� �g\���y����=�,������z�L��++9�NeegW�֖\��PPV�� ²��^�N=z���˫羘�@������e���a��C���i_��S�¡ϯH�NN�Gbb����ܛ��f�p 9�y�tɽ���̅��Jo�ULF��܋�~�x$�H��L"���z\C��P���o	)(`Ln�^�q��8X��"��'�V�	(Zv�@O	yxx�2�4n����� U_Qk8�Ξ�s�r���R�Y�a������X;���U���ο�����Qc�Vr�O���������}��WTT$�� j�MiY����ɿ������~�{52�$k�*&��Ʒ��rZ��R+fY�J=�d'���K�~���)��aݷ��N1���!x*�xZ)�NjW^���A�Z)�Gz�`u�)������3��~t��Y�"�X�g��̏4A�y��z?P�a�4�FT��E,�����43������|A��M��<X��pEʍ�+2�_ T9gx&�w�8��0P������i.X�� @ۼn/B��j�(�J�Brg9{{v 0��))�:��%�MM`0xx��������� �Cv?zu����hE��i��.;>;��+?a&��l�҇��k��;��Ƿ�C0?��l�{U}wH�Xf�r�����톣����I����fa���TU�E�x�|�II-���F�5��\�����$H��m���b `+��t�1���33}���l�^����4xaE�������l�'!f�]]��q���φ6´G����y,���2QL(���m���iЋ�
��yy<�,9���ю��|���DG�q.�����ڟ����2�z�5�Ji��H�:��������Ӎ)y������	g{4?%N��8�������lHE�n0ha
�O{VG[�����T���c�iַ����a/��O��p���u�|� �O�+����C�Ԝ�=���y���##�?����sȔK���ָ�l]����Y�}fzz�?BZ$�߹Пi#�C�o���9+�b9a��A���� &#ž	�
�W54TVWO���&<4Sk��mX ҁY���YU�^m>�Y��c߼];8�G2��m �@�P��]o�������ssr*˅D��)�"��+9��NO�8e������DP�З	�����9���?����m/|���qu��(�y�ɮ*���SQ��Rt1�%|*Ɲǅ�\�@:'��K3,��"ǘ
]^!B���ѷpc;΢�-�ڊ�ЅU�@�8�r���;[����2�:*?�"d͗�qԛ�a�IH��ma4���h5 �N�l�@�iEr�)�n��vܲ5�Wqr{j@�JW#4�V薝���R�{��wKaƂ�E4ܬ(z�����of&�\_�%�:���n��g�����ܠ�wK��)����;���]��gyS��k��aH�g�p�˞�����ሪx&��-����666&nnu�:���.v�YW~/[ʧ��6�6���9s$A4��U�..�c�5ٹwxP���b���";&x�+����<%,`�ƍ�WUꙔ�==S�B�~\�l'཭��5$K�����"~�+���x��h���ߚLsD�2}A��6�N�_"���zɨ�#˲��J=gdb��u�}� ���N��_j�*���P�Ӫ�Y����6V�4���{�
Y������ldIZz�s���5Z)��0�D��n��]M�E�ːq�:�挚�(�QYm�i����.*�WQ��eN�N��׻J��ǐ���z�ZF�1I4 d��/���}��9S̓�C<��)�I#���K4j�}�'�>�3�3 w�lo�;L��YHT�E�̏�F�vCҁY�3ne�>3�6�g_��kұ+o���K��w�F�^�ҧQ�&Bx�����������ƭ���
���$�)P�DO�[�#=ې�*%2���郉;������9�$����ӌo�n�����W8���&ja��=����k $U�
����sPWI���2�K�(	V~�<��:�F��B�`��!��ApUӲ����b�n#_���5�q���wyFy<67��A�ڸ�a�|B��H��=�u;Qt�(�-l�xb�֜�p���P����g�����7jAޕ�o�}�����.�o�j2�z�&4D�;a�Ôby��p�Y������j��t��2��0wQ�e Lڞ�Q��z��>+q� zJnUѯ�^(�?��i�hZ��Ϳ�J`+�K���� �6�;o�7Im�'L�l��K��}�Effw޻z=%Y�Ԝ�m_�|�šW<�U�D '\�z5)_*_Fӝ�r�.�r�T�@(u�_O}2��������.<ݞ\={J��.�ޟG���蚜�Ǔ-�#�]��ě�-an`�Z�EA��	�9�ɾl0������n �nCɩ�a�>��b�,n\̓�k��{����������D����������b*�a4��,S����9�s��l��h崬��q=���`K�-Q{kX�A�K�ы�n��d�'V��'������B���kv���I˾#���_M&0rj���q~��tk�:X�:�#e����8�8��C	*�9kR5%e�3�x��X�Q8zx��]O!K�w|�����̀�Kq1_1Rp�7zA�����4\��o4�A\#T_�x��mn��V��'3�pdV�h��z<�q$��M1�����02t~~�W�J�;�s}��8�|�@F$�'Fl�p鸧�h����X��ڇ�b���945AT݉�mԁ��Rb6VT�����μ�=x�L[+������nAO����o��6q��'�	+'��}��Z�#���s��]uF�1oݝ����߮3[	w�w'�7��X�����~���)M���L5�d�/�+�ͥ�LaJ���d�K�n� S�~_#�<�GW��B�ѽ�JS���-��e}�N��!詑 3a(n���O�ڛ�����c%��Y�+Nd��~�a��5���l�.\�J�#�����)AG���u�t�	�v�WY��r�I���6�f����q~��Ϥ�0�vV=����Y����Բ9-u<;�C�Y��Y��[ۇml�Y���)�����x)k�H�ZC�k����[u�!�4=v��}f]u�� 5TG�^c�y���u�o�����t�4�Fk��؞T��#�D�+�hu��Z-��S;��O1��Oӄ��}�Jw��U�v?t�6ڇ�{�}j�g����02
�AGE+�kېS+[W:�e�O�^�<�F6�]��SS��]#66
�6������vL�C��LW�a����BKlݧ/�7<~�<c�>XĩR|��#}���ݫ�=7��8��d��4��Du��$l���5Sk�x��qv��Ffq'��X�p��\������ޝ0'A�A4�,		I�3;�*Y�1�ݵ�wo�ީ�y��C���tAqtU9Y��ɓ_���˳>��DaUD�g��*,�mɰ�irqE��:L���0:m>��4Ϸ����F1H�j�+Ļ�\��� �9��+n(qrbPTtl�FZ:��_'�>B����M[��z�BddķH�~�r�coQ=�[�����>9˞�����)�xZ#*�1rm?��B���"\i��B?�,��[���D�	����l�����E3��w�W��syH��A���R1���ݔ;�@�1�0��pMTb�ܿ-���|��2�����n���R� �g���ހ�c(C�Ӑ>��*юc�2@�!���~^��Uz�-`��R+�+*־��鼏i9��}R��[�}]n$�+��w��E�T�:N�Y3��[~>�t͏ f�@�"�x�}=���Ѷ���������6��J �oK�E[��2��ڿ��l��c-��� ����J 9�}v�ڻ�dB@�];��v�%�y��~�(�o9�V��=]�YF:���a�_
1�[GgKތKd!R����C<�3i:y��7ۛ��s����k��s�ٴ���bݩD%��/T拢D��#8s|������O���ڽ�ŏ��j��c:Z.�B�*��:o��Y{�h�ЖdSާF"~�/*���VH|�����k�Ɩ8�6nr��e��K�ɘe:��$��"ЗH��.����7��v�;��^��a4U�K���Eg�`����x��M�8�R�xJ�gi�_�UmT��΂�����0��<ew��0e��d��]�f�)���Hܓ��Ae[`�z��e��
y��cY�bv���Aȁ�[����Y�V���b�ee��E�I��NaWIt3j[��bRQ#55�Ϫ�b08E�YP�j'�"w:~�Y�[��))iLl,����He�0 f���N]gV�7[�5,OƮ�r\n+N����G�R�MW�y�i��_#〙�<HW2=����a�~�w>�C��!��_:�h��F���*�����ؚ$R���IB�i�v����<ם�M��u��>�0[�}a�_�8��J�S��@�?ꈂ���e�
����7����U�,�l��T�E��ӭ�����=�!���L7���B�	�0��տ���FF��?�������!����*�����������N�wXDpxk�Y�6<]HӡZF�*�j8CDa�5��=�?�u�����u�5e%���W0n�k|��X46l �v�Ŷ�=8d|j�7��ͽ��I�XM�:��0D�k~%r�c��3�ی��[eGC�Ez8��Bb��K�Lد��3!�6�'?_0[Zܶ�r��]�y�Tڎ:�/71��њ�+����}�՞.�E@)�.�߸�@��!�[[[�D$����4Y���ˆJP[R��� ʸ��1�������7�W�F�Cc�W�bg(Es��[؝�ï]{'Fo��n՛T�۳q�%RvqL�����O�~�:4�?X�n�~��zx�.��B#I��J�0��|��IXa���'#���$�WS\k���Q{��	��X���-�d�j��r�Oy@I[G(��.)�S!���ΉcY�S�W���~��m08��w����lla��%[X����8o�VQ�t�'���z'gR����3!��,�kI�YYsvޭD<�S?ǜ��Ț��i[�G�^@�����N���Y�B�:D�;3����������}K$&�����:�7522�q�v&��j���ڢ�K!�܊I��$�4@F�l�I=���i��^D���_Cd~ڶ�0L��GW��m�4��jg�ȷ��������!K���w4��у9s������=GDu/�jDB���Yy��1G�����7�I�΁ژ�N�u�b�Tp�̧roy��:�X�9�J�)[����`���r��5�7�#�"��J|qrr"C��zNpnL����@~�����������H�1�?	�/婣:kC~9���	U�F�:|{ K�9�o��ڳT�&�p�Ou����`�_go��Cܻ�]s���V�ӟ��@�r\:��UV�=����xgH*����r���~�W�s�w3,�_������[�_���E��@�:�
��d��<��<�y`��zi��}	�I�H������;8�ǫH組^Z&_�$��1]�uKQ��7�C*��|rr�<��K�N1"�Q���n�B�1N������ οVb/c� �ʛ�C�2�}���W��CS��M�[����ۮI�i��CJ%ͳ���o��l�k�W9�X��̨2.����.z��J�盅|�Q��͚�U���#��0�t�NGq��f� ��������>�F���o�6��Rܫ��7�K/Ȋ<���/���B��'ㄽ~B�h�]��������b���d�	��/����g�'����rg��T�����KEO��L� �r$��>��y�i�{�������p4�pg�UWS ɷ�a�7E���D �[���:V�טtث���p�Ek��q @�hJ�#u?��gg��o�z0�%Y�%���9P\�\�I�m4�W{�)��S��������k�-���\Yנ�][��4��V��G���ھ���%уx�N�P�aA��b{�b�Q���6��<�����$ynR��)��C�X�ֶ��� h��|��=nir!��7q	�籈,�F� K��>{��s�y8��_Iz[�[lW��[��T��)���/�N�'s�65�#��9��<0��)�;4�H�o����-��鹲� K3ʅ���	�!�Smw	�b��CN!�[u�%�3��٪/��BoFn��z�{�/�<�2�_44H�	�z��Y�E�^�%�V6,��K�6X8Q6l�����ct��y���ț���
{�0y���Y�1��y*<v?���k|��|Q˧t��>���S�����<T�Z|>;����w(ޓ�ƜG-��w�C�GEǋ9�S�.���rֆW)��i7�NչV�*(�`s��֗�f�������I��C��2S��=i���^�����mT߸�����M�7l���|����ai�z��YȥA�J���E�TFg8��C�Z�L�P����}���[���6����]�0t��%��57�s����Hk�m<�=q�DL�Z�W����������So9g0Dv\\H�9���~��)K[6�)ЬA�d�s���p����Q%<Lo�%�V/G~��u˲��G+~87�GU� Ro��#�}�Ԍ��������)�GR2�$���e,R��ajA�s������ЎH.��*Phf�B;����/~�>ho}/`M���@P�:�Y_����ϵ��M��d!aI�7pm����\[�@7V;�ao��Y�XX���O�W>���P<	\u��mVR�7��I���ϭW}�R��X�Ğ��tx�Vs�E�sA������@_g�,&ە���7*��mS�L`� �L������Q,�ZΗ���g���U;~x[�`�K�����j�*���z��U����ؑR*�R��p}�%��R�����/B��׬������/�y���Յt޽����R�ٌᬫ���%�����u[��A�P���,�gi��hk�+X��L���ߪr�<����} �21Y�5�UH�~Rɩ��� z��&=�N�A�M�W<g�w�{e33�F)]�g��(�Mp�$?��1�� ��u��?/���OGZ[�n$��7D���!�s��Q��)
�8�H"C�/����ݙ3�i��u�m�+��WF���	��,�\�J�J�Zw+�J�r0|���?��D�!jM��VeN�,����L�������'�s�n'�:ưr|oy����:;�ݏ�H�B��M�"��"P��d����g��힓��s�����w��W,/4�c�\�>���oo�ԡW����pQ���Ӧ�/���Wmm�@��nzON[=~d^q�[��)ok���g�RN��&O�U%���^�!�}��U�&@
&��EwSRS�4Ǵ49-Ku_��33c�ӏ���0ɳe�$f&���wH���~{�:�Ɗu,jk�z{�U�N��\A���*�^�K2���#�_�z"�.�o*�gY+��q96�R����L�Cj�OP�,�0{ �NL<��o���~S�M��[-6j����T�f����TÀ�u ����C7'�e�'O�>/Z����n�+W�7�v�ҳu�$���oHb��9�{��\'W�#]P~�1�oxz��!���@[T%A�Y�>�K����+ױ�,���k�k
�t��@ ~q�J�@�yN��e���ikv6*�6A*1�Ǩ�6/�WV&bR�rj�GN)�y_�/�������?zki?豖���)Y�$%*Pa��k'Y���D5	�&�&Y�'Y^�'.0X$f~���@xT�ZrS�x���"P/"Q�[Ιw.<�v�@/K�9���F����Q������93E+F2\c�����2�6�>�%�W���Qx���D����άz0k����ůؘ�sP_��ҝ#�;]oKQ__�
'�|�:.1��VAY�Y+?��%�t�:�#�r����ݑ����@�Q�op���=��o}f^�[�B��f��ؐ���P�=��O�w� ��wWY�a�2ғ�7��YU����`�Q�ZԷ75 	�U��]R,[�K��(l5^�҉�% ]��!��}Nm_�����J&GF�ݧ�����>�:�œ�� yI/~�*))�!�cd����T��r0�Ľ�LG h6��P������� P�������y����C� J4
��N����щm�l�ePx��t �0�ְy,d��ZvJ���('\�R�f�~�miH��X���$8�{�^۪�}�y@~����g�x�a>$|�&/gkm݉h{8�b�^G&t,$�}�@��	o���_B�BE/7 ��u�2���v�<�6��z���TH�%%~�VCFF�SM@��T�>���:{���Z��Ti>)]0qrz:�˿"3T��t�j���I7�oIL�.���</��+�؋TJ�?1�G���/�=?|HD������X'�����kk��I�OW��MOO�-i�Ju�o+Z���qы���eF�To�f�x{�ǬQQI����7�%%�$��� 2�SXY��W ���.���+�7�����}QB3��,�q|o�4�C�UEkuu5&&fdz�a������ie�ew��WG���z��@�O"e��zW�;BѸ�1a� �󙽽�-ݸ�,���`�~��'A��gD��K�g�{�S�B�#�1�צ��y��^�o�8?'��XT�FFF�~��X)�{UU�J�TԷ$bx����R�/��NK�9����/����8@;\�_w W��>3?�9�+���)�ßG~F����2tU@�֜���B��d�7�}fc�U*��ִ�e}`,12WHŋ��T;���{tu����'=y��i�<Q��;ט󗖖�޿�1>?_Q�%S��Z�YKgM�˿?��#�x�.��)���:;����ʛ(4E������� �|������j���SV;:??��*^t ���@=�Z����Bn���D�qBV�˄�R/q�jtt4+��Zl�=��w��N�� �d�;B �&�P4�z����-�+d�����/�JMR��ҽ���H/�j�ht���ں�J^:jzpPA	�����r�u
嘝$Q�ͣ/X�Ց�<l�s>�j))))��%`��#/���NG&�� ����b׀�����Uԁ]�xiFDD�F����15���{rv��-�N�N�e�	=���	��^̕1��t��u���@���R Ua�r��?�/>JݖR�Ft|�|*�d4zJ+���*���_LlF��	��4�Yǖ�,�۾��k��������.
5]8���'Ǉ0vRN��롹ۋ���b(u ��w;����M2̏}NCa/�5��9shH�V��m���sf55[�|g�I����:���JP��"�X��P��%����}3��
��I��(-kj�f7���^�<;���K6�?S�~�&���NU���s��#!tԮ�òQR����A�P��Y鑗� �/3H%��!�m0�ϴ!ad�+���<T֔�n�W%��z�o��>���:���*���g�~�A�p�Z)��F 6�|�h9���cD�W���؇U�Ji�򛞊��Y�F�X�GEkk��+x�dpzz�<EB���X�L����"	�f]!�V_0*̜��s<r(r6�`Dy<��}��ψ|>��#ڵl���08���_��񫃳o���҆���;shM��ᓧm�Eq�f�b.r���-@2� o���Sy�9G��o��\�p��3{��D��!�5Ԕ���`�%�C8g���@5��i�����*/�~����&U�����S;��]tK�ۨ�q\ٝ�z���]���K�t� �5��b��v�M���Qz,�f����%�WOH��_^
�kf ��Pl3���F���7�XZ2���gm[4 �8g�夥�UE��hпO*J7�JD����R��``6�T�y���?q���E�u��:�����4g���7������YT���^���"���)�`{xMN���I����u@`)q�J��<���Yww���.@�$�7�W�2�O�Z�!1����tW��ǣQG�{��,������������V]���D�˘>�+�`*XV�k�,������L{	/��������c>����͜�%�������v���ӟ6]>������Y�U����YNww���Tߟe�O�;�W�Ʉt��?�8�<<֨W���B�(L�<�o��<Ox5�9X��b��5���K�4�cR�k�Γ����)R|�������(�ہ�)�:
۞ɛ�wI�����j�ڷ7��m��\:S_��+l?�A�5n��C���{z>�����C����$��{j�R�HP�(��z���w���B�%����Iyci��:���p�ʤz��6�J�AŨW ��($��Ȧ�[~��>@�=q�|/-k(QfS��ז��qPsqO��`����OB�"����M����<��b2%ݦU�:���q.��?'#ݟeL*U�O���ָ�Y�TQ>�+?)�F����U\� �K%�b���*���*�&��O7V�^�X��S4������
%���Z��Gv1qq&��	��j,ɵHlt?qC�	�\��A���U�G� ���)q�::�I"	ʏ����j��<����"���D阒������袻]<ĉ�)Áv���i����	z"m�hh{{����9]|��/Ͻ�����&O���LH �Ԕ!����J������=�9�D���!vs�� �JHH�g��V��`*ZZs??�S�ǁF�0T�N ���Wk��GJs����)� Lal�zhny1]gM*&&�ݞӻ�n��l�a�G��KHHN8����Y��5+Z��>[j�O�݄���d�;-6ؚC�He�F�_b>n_���j�_���0��C�}�'>>>%%%Y� =gea���VUu\=P�%+:�	��ϫ'�������֊����[���� <�e�`��3f7� 7����ҞQ�n��$�k'�H�0S�r
ʺ�"k���`x�F3ob- ���
����O~;ݨ����x1eyy��ho��g�OGFG;;:�"�M>E{0&lڌ;�v�q�ܗ�X�{��k�6��a�G���
�6E���WpPl/]G݋��w:j�rsP~;6���3��'��� <�:���\Z�r>��� ���YO��kq�ڣ�pc+n@Z2��3����ᅟ��������+���*=�
�w�j����e�7��}{�
�lO�#WHb�����f������	{ʐ@g�A��<����1qB�( ��g��ܬl��!�5sn*��ml����-���L�pm�W�[�4e>�~�݋c�S�rCҦ�i��E�؞<��K.MD6M�y��HL�k�ѥw)7��lB�D�"��as{s����TQ�}��V;h){�:@�H[�kW��t�뿄�p�W���r�1�.q�T{|V�g� ���@j�}�3����B �	��s��;������a�����4�,=&ZZaoEc~���ؠ02���d��{g��S��}�o��O�8�K���EL3�Z�BIde�gon����,���Zy.r,鸓Dt�I}�þ0�gZH���_oB���~�nn=֏�	e9^}�
�}������!������9@�lV��d�_�mU��������\���x	�Kz���LJY���ܘ���$�ǫ)��=�D�8m-6r&���l�����ߟ����([A���"��YA��F����sv�V�o���;N|0j��.D�ՔQ��>Ԟ��+-���):�oBL��Z�$K��	�vR]ߓ�n�����R��lll�&$|Π^�&�sT��% @����|ck�ـ��0&[��W�%ɨ���?_	e��!����?z'뮂=����-WA
��ӡV�Q<
�Qg�f��#^/����ؿ7�F�R�ɷ�A��ޟ�jkS)e	�kq	*Y3}����#Z�L,[�5�#��ψ�$�j��_�%5d̐1�v���t��f�F��ϋ���%P�ɻ��zrt�8r�ׅ6���}~"��(����,��ۓ�^� ]�7I����Bvw��i�NJ�2�K::�x�|IY����7�_�F[�~�Ɲq`F��%��e���ք�O�sy�}����_�ė�S�$|�f9�-��-�K����vrru�����[��#��v���֎�B���t
׳���:�<`#_��KLR	̥V5%tL@~�h7�x���>�6Oxsy3��b�{������[�C���h,,��߲��� ��%���� �؛�S���j�jo<�4��]=�]�%;:;�0���ڛ�����V��a��C��1շïn���F:��`(���-���Y�f�����kJ|�o���&o޽7ɭ`0R�0��wr�'��xm��4c��.��l���&K}��/��`:h�m��'�������(%k�ɬY����M�>;_w6z�Z(��96zL�XHI�2�����]����ֱ����9�E'�O�P����!���W�gQ�#[~�cBFA��u��54l����muL��e�hY5�n�|�i6,�{g�������8<z��4|05�.���BoXOI����b�{�xu��95�&Dg��n��R�������ӊr��!��ER9��W��x�R;_��>6��ZR��7�,�gw���֊�O�{w��m��+E6[�N��د���gs�<1��^+ll�XPxaX��<YU��S��f��w�d�lu?~��?@��+(c�~1v$��ۛ������SS�|Ţ���8���J~�6�ر@ʨ:p�c?G9���aZ������^������A�!�zM9�X��Ba�gQ*�]]3���$c?
>�V��=K��?tB�|ofF������2~�����:wv�م�=�ҧ�%
�K�0\�O+Z���y#�p���yїQ�:V�ٵ�墩b��k<"�����M���|	L>���W_1�i�L�~�xsx����GxI�<!J���CKO��/�О	So�bn�?���+��}�ghI�n�S�A)AZiA����[R��f�n��n�{ȁ�9���{���	��Z�8���}]��g�B�;��!�9�0��K3W��u(�0� �a|��D� �Z<B��߳�z�A�J��2z��X�����l.�ʷ��+��x���vZҧ�!�����J�9	�x��.~>Ps�hj�%t�C�6<(h����O_W �+՟�q��Қ�����+DՆL
T�	�de 0��G߻��3v�:g=1�TH�5)�J�ц+�~q��_+�� ����i��cס���P>�k޴��p�A=�ް;�=�7��ġ��AL�regI�p�ճ2'::�r?���T%�:;<�!󲪪t_�C�@�����@o݇�������p�@�͑�Xd����O���FS�w�\�ƚ�˸iB��3e����|�Ut|��ʕ��m��>W�0j9�����j�����,��'C���eCs�t�t�((�8ዙi����V˲!��D럧�>lQ�E�1�3�d�g����J�RQ�D᧚&�N����򜛛���e�US���,-M$t\��$Һq�\|.r�:��ް�>�t=��]N��['�6%���[x��s�5�%K�o!�~la||�7�S/�1��Lq����d������Bz��� ����@~�KtK����ed���{w��`b�C��S	��A{ TS�(>H�kK6تf�mv�z�����C ��;�{AC�,���b/~���V&��5�����U0W�c7�--�r�0�X��x�k3L5%$.x3�'J`b�6��yJ�j��s�h U��(�"���{/�Ze�4�秔�G[n5;CT��y��bBEe������
rl�	\��A��tN$�u�	h6�x�Sx�'۽)�
y��{ ��_� �������T�W��*�I]� �(��ϳ+--�]�R�CD�/��-.X�ӂ��5A/�kP�1��ǫ�E�
������a�lfE�َ���{^}ɭ��+*"u:���	��M�%�+Y� �Ix�Dż���]Jꇱ'D8��TLL��@4���l����|��P!��o!"3�t�κf\��C|V�36]/Q�+�:~m�q��*\|�5zt'6{���ށ��U�DE݉�LE�DZQ��*/���Ej�:�Q����6�~�4�{t𸤷Jp�{�|v������������18Z>��8V@JF�WTNd� G��v�F���	���V���f�vs�f���]_�Ќڝ����u��c����0"���U�TWp�d/%b��l!�;C}��׍Z�J��X'�$B��R��{�+��c)�_���4�d����� |bͰz��l�RBB�k�k"d'���ݸ�Yǋ��\��j��0U4���Ơx5��S�٘����崖�Z�?^�~����ϯ��#�(�89��8�u�vU3��g����D}��k?��Pm���d|����xh8ᗞ(C��1���Hǁ]��c��疸w���"�g }�Ke�9��7��	��|�]on'�"�f�������%�x�tph���� {&a/�hcv�3!}��X�~���t���������C�dہpL�Ï�����4�NL999�}$��x˶a���O���	{B�L����P�����%c�fkK%�1ﵓ;��1��ş��0��6����r��`�[w��Pg���ml��vww�����ޛ�>#ľ�*�I�:�Y\����/������ba���@�x��Y���'\���j3�N&�`Ee��v��Hh�|�m~�H��mq=�/�(�[�l;��M9���9�t��ۭ�qr1*881���(_Z�f���t��t�o)�V�z��1�p�$�O9.�޹�'���a./B�oPÞ:�w�� ��h�(Ҷ�V��i�m���ydGq�d�K���!֠��"d���n����,�h_���62��}�)�a%���@��qP^T\,8���UECc�f������r�q|h�Q��z��ԏ���z����X��J��lD�6C����&D���T��X�ءqۼ�K������>�"�Ӵ`�TTTB##��mL�ssr!�g
���6�\̀=F�Z�S���E�|$.;/R}t~n�TF�V=�w�Wϳ묔.��ai�},�~+�i�}.�ש��D�1ݤY�_��:$Z��t���N�Hd�Nb��x��w��R�)<�����;����W����{�v�R�H۶���҄�1�?�"����Yn)�m�c|��S����TgK�ŏ*:� �mtZX��Ǡ�%L-:I3>��\��Ӏ�idК�We+��烃�NGD踔���J_!I�V~��q�Z2������m�{e\��S���"���2Tb䔕��q��������U�Ab�6�_J����KQ�9���i�de
9�e�OȰ�"��0�
��η�������
Ty�E��=�A�ձ�y8ݷ���]���SBחHPr�����P��,� ?~�Z!!��o��+)�,)2��n6 A��(�M�B|G#�����#��zڢ��+RR+Q��w&T8'D�K���1g��`��G�$x�\�������M��$�|����A�=!�+�'}��إ��q�Y0 sd�Azߨ�=_D6�3!���k�A�u��0{H�60�S��f�`����_���	ˈvpq?h��izw�QiZ<��7��8��gS��9EA��;'@b��fC��@�㡀l���gT�UU}�Ջ��KYQ�3F��A3��L�R��o���9���^~b# ����T�\�Ea���Uf���-d��v5���S[2��{�ȿ�%X�v����w15�jm���L����b H0����1� X\E5�����]Z:�ײ~ԥց+%��2� ڢ����,�g���
`��PMȸ�ͯ��Oɟ��������x�Ƙ;���*/��M`�'2�õ/�`*y���o%A������&�P?���3S7i;/�\��* ��gtA���ߺ�^?��fG�;�Tr`����z�{�l�\�A��p�����fç�c?HVؿt��>�g�^�ɘ�G�}�5��?
$M�6�ь�la0ˊ]R�UO�XȁT���(��:e�����HP���t�W�+D���b>~��[йXd귲��m�15�jq /��uqA��4*2t�
��}��]ѡ�c�����U���|BB��N�-ˈ��=N�3�G��S~�"���"�[6˿e��/��vr�T�P�r�����������d���� �t���z��d'ɮw����J?�T���%���Vo<k�gץe,@����#��pQlԿ�H5�3�b�Qg%�Gq!B�p�o��ܩr�ıhoP��<$�O@%�E���S	���uio�W����z.���ޥD���S�G��]t�h���!����3k�ہ��Z���~�,״o�W�;<��t�����
P��/�0������y�n�4U|4Ee$s4,gb��U �{4JvgqM]�{{M̹�%
�<���N:�Q���%e��{Wg*��4yY���B��:��=��-��]�!�4t�G�e����� �̋���b��v�+��X�N��j�B�j��#9Mq�M�U@�NK+G��?>�S�0ꋰbNR��IW�2KB�ӏ|�i
�HV#M�+��,,��{'�c��bwB��m��
L����Hne;����qI��By���~<�~}���h��v�����̤���ĻĬ&c���F+!��m����Ql^ggh�����]�/c�9tO	r�@}}&�������f�V}Ԛ���'�P��߄�}�#y���=,0�B�׺_t桷�\�y�IKS�����n6��uJ����������ÛN?�N"��j�7?�ʫm�R�hQ�嬕�)�$s��MY��ts|�U���Ī:�>����"DJ��U��x��l{}O����p��'"(�#����^��j��N[��:9����zuT��x���*,:�-!��Ŷ�ʴ�/�!�S�~�@Z��#q����
h����������`,M�8J�&��,�1�Wr.`(`�Β��T5n!9�O��꿨@���/��|���_[��v����`>�r�㒭o�<*�N���"!/�޷���Rup�WNI#�ȱAy���@G�2�%�:�]M���\;H�d��+]HZ�^�� Z��C�:m*���4L��5�D0Sd�>����&�B5��y�5�,�cӳD3)F�Ƞq��%w��޺v%؂��.�^�2�,#ߋf���-�X���_[���y.ق-��ޫ��H����:�o��w��Z5T���U괼}$�A�0�ձに,�c������6�X�J��%��,�,8-&�o��Y�~H{��)�%eUQj	GΙ��.�~N����n,�NB������$�%��Ǭ%E�Z	�cM�>k�S���w\:���2<��7�-lؐjȿ�p��d�n��9���;�Q��Ъ�u	,L�<��s�>C���g�n(�hd�����λ��W^J���_��>�R>�d�wa �"�ZG�Ү�A���c�G"��r��i���2#2�2\{0+�Zˊ+w�Z8EQ8/����K�@�K���N\�^����/����x&&&?�����01�j�R� \�4��2�YI?ϮX>��Vm��kl����_�).�YO�b[z�Z��W�T�U�f]wR�0^A�1�f��,�)����c?��[q������_f�4 1�����녖�9�A"r)������}P�؎���o/ &���;�]���0��}����__O[��&��!��ߎ8#�]�?�'�1�i�@u�����3��'��`�3^�+�=�oib�ԟq�|C:�ee��l����46�m|��B�G3yY�����D�1+��PWd��zٍ��-qd�����6���;�����/�L����������L��5��9�3}ٟs@A���Q������޵���~[�s%,�����4��5L�TT���KTTU7�A�/oDL�?��J��=�p�i��{(3:.�t����v�zJ�̦^�j��PcQ�"G'����߈��Q٬�߂7Ub#S�a����x<�a��2U���A_.'���1o'�zTa'�UU?�d���ϫlĠ�$�a�<mۀ?HN���1`�3/oB��'ѕ���~���Ryq���(�斴�im%�)�D�Q�j�+��Y̠[{' vLۤY
l!58]zY�^�A1��+~�ݴ����{���Mϳ�]W]��^��PM�2�V
^����E=��8��-�-"$z�� K����ĥ�R���}8��$�5_������=+VQ�T��s��b@���fy$�Ң���4u�ZΡ���a��N��\�s�p�~�sUf�'�����ޏ�G�ܹ��pX��ӆ m%�)rWȒ��L��5�v��;g_��Kd�<PR?k�ŹϋV���G^�D�}wq�A� #���9��VJ����`?ZГ'#l�Nug�?hG;���v��jm��hȆ���+э��@��)Z������M��z�9��
��r����)L!챇�x�rK?��xb��z2�82��Y:�vȱQ4�WD�x�`fs}G\&>p[K��z����P�uE��;]��@�x��3ug2�p�_�����+��]��1�v4�?2����ɶ�Wu�Mz�.a8ho^b�5�F��)�pR#8c�Qx/�s�_b�9g��G����k츼	���x�t2#�q���qE��J5���쎇mn�B��T����_������e�4��74=�2ͬfmVN�����b5�a�����֬�<E�Ƙq��E�*�ﻠ��0~$������Lg�F��KJ�����(v�Fu�ev��.������l�v�Sg�fw�����'�W���a�Q�j ���.�xO�a���fa�u�#�����L,��4QsM"d�fS8�ٞi9thed�]d�B�Qr��F�7#?�寯k��&���s҆���,��"�\h�1�>­9�b��{�����ղĭ�ݥ�n.%����5�@����vnC���{��� @��+p�4�z��;�A�l�P߻VH<����¦��T�t��F�F	�OF�˙�?ؗ����J>��%��Tl���?�YoW4A��V;!�CfԿ�X���s\����}�5i!�4��s+���CL���Bez�U�ko7[�*v��9�zX�Hk9_,��XgNF�C�팯�h+�n��?&�(��76N�ԑ��+�S�^��fm�M�,d2�g��E[~�#X��O�� ;I��Kj1V̢&��h\U!�C*Fk�2<��3��M�2MjAY\�;�/����L&=hxȟ�둭Hм^7nk1�f�)b�����O�@��8����K��'Y}��Hs��

�ŘU�n	��lB�z��}�$DL^����""��ozaR����X�w�N���`m�c�x��,��S9
)I[�cZ;�LPm{��z��HߡS+Y�����ޱ��ْ���~����/�̻�:�]w�v�w&o淭�:��w��пX�0{0l@���3?�}��z.��5l��$����K���#�H�1}[���,��>��`"K��R5��4��Zsº��6oա��1��BR�����&���/qx� ��.��)��RBL8���LW�E/v���Ԗ���S�>FE,JeЛj��`a�N���$��F�k�����P�_���Hb�0(��}��de��@ph���&4 ���"�;?K+��B���~6�Jj��1u�:�.�oV�kL�����H�n�!�B>�x���9_��8]9�	��،�nc��h��M��0��iV�����ڕ�?�����)�~���Q��k6>L�����������ޙ*��t�L� �5�K$'�1V�/c�9���֟���wXdNE�~�d�n|I�1ٱy�D> �N�oo����:�H.����Ҋ��d�;�,� �Yvd���X�2r�����V8D�{K8=��s�^E�ɼ�'S���D 2t�;�7���G *�P�n'yhF+qҐmyo_[3��o�&��$.B��Z�B@�M�h+O"� ��d��s/h��:��W%�1Z ̷�i��f-���Ų�.N*nr��O�� n��Vu��hVN� �j����A������\���S�0���"a�	U6NO��������Ǆx��w��������7&��E���[ �.=4���GƲ�����p�5J��Ҽ(l��������1�A%��Q��X�^,��9����aoТ��U��%��Z�A���_�F�t�#t;A���F����鿦��5���W<���^M+��ܩsi��;Tp�Ao�q���5]�b��E'�
!C>�ο�D����p�l��F�]��KQ��&4�i� �g!���L���F{J�A�n��,,��6UH����]p:#@I�k��@�&��a��X�Hj��;bZ��N�� )9��ߢ��w�4���#4T��_��X��k� C?���0���������	�h�?���ɠ�Y.x�$h���&�"�ҟ_>�&��

Ҙk�ă]mwU�Q���a��'��Q�; pCB��F��(��>���3��^K}W��e�ϯ��'��\����mP@Y��h;#���ǔ֋IA��6�{���s�h��zl��3l^�g�w	�Oô���3��mD,Q�x^��x)��������m��8���H.Mh����2����_�GbG��#hO̰���".z�B$�b��vQH��t�4 F�ydg3"��t�����O�s���;�A77���*��T"5g�G}0}jr��˽x���R�«@��ߺ�2�Knh����UoסMdt�ь5%��+�#vPѽ�3A��G��(���Y����x�X��N�ȥ%�^���������S~�,��|�~5"��х.���/�L����gCq��e����K>A'&���>�̣>�}T6��~�K1S��D7��Gt~hH�M��Nw�D����)P���QE���z�Q[�\�nː��Ñ�^�sQY��4Z���r�Y�.r|��a�Ą6!�f�u�s!!r����[v}/�d�3L������
�:�a����E�O_�ƈ��+#�k�0#��y���sn�gaaz\��$��[�^g}�7k�L�:$zSd4>n��J�й����A�\.�����K��:���;���&�(�:
��7j��Q�O)(�@򊑽�����ޫo���~8�n���l��<�淡{JB(7.#i9l����̇������<��:$ee��<փN�/��v:��4�P��2�0��/�ᯌ�o�t�5�|`���) P�����c�͘ ��QBO�܍Ү����GkkR#㞱vo^���PncU*�ga0K=7g�𻾹�=�Zhi"7�s<��Sx�E�q�K��r�F`�q�ih��~��	�:=�,�?5��=8`x�|��1��H�ݝ��;����CC�O�}�ɮ�&b3b�yX�磫p~�d��h��A��R�V�CM�Ws��T=:v6g{�0���Ka�0ו[�f������]i���u��#3M�]V6�
��������f��aE��~�dvI�D�O(lw����Q4�x�<�����DЁ������eP>��ǂ��q�>\���?^�Jt��|y�W�ѡw32�0��O�����t�����nha���#,�����@��IJS�>�W�9wз��In�ސ�_ŧw^���0Ù2�h���4p���1b�5��1Fۿsݮ��n�Ȯ�1rXO�����F�v�O��'�o&�$�>��2��R�j��zD���@�.FĽ��}yyL�7�G�<;� (! ��Q�y������V��;������;`=��Sw�Q�2c�� ���d�T�%U���jI��/���EC^a�S7���ل��U
9���+�]L������n�K\��~$�$�B2u�|�IT�����}(F�������n���o�=O�N�.F�p�c�pz��iB�B�o�ȧ�Ĉ�ך=Θ�08�%(��sz���o�Pp��xLM}��|܊�X�;��\v�|�����OS��������l{Gk=����~��`o~f�k}_o��#�������oQAy��1=|�^ٻ���		� ����%�z�$���g:�����Q\�s��2�W�7���7������g@3z��m/�s
�����ۨD�M��Ϯ�%ӣ�?*�ЄM�o$˓T����&��
��1���}Y���V��ù����b��ч��d�ч	�k���$T6ݍz��#d�Ǉ�U�	���r;#�io���<<s����I�G\0@���9����A!y2F���en#�� GI���ۿ>��?2M>�P�莁y����KO z���,�� �f�%Dk��t^/#Mz����BA���oKn��H	�бAY,���F]&]�	�
\V3�]���㹏j��(cĮ��ud@�Si��%��#݆�͐3Oow��?�|�����"ɧ�?�̒�ޟ��a��|]�c��-�F,�=���$�\9�t�����S��n���L=eJd��~�Q�O&�݃�tYgH�k�Q�7��Z!���j�u���h�����we��p���1�SP�d�u�}"�T���)l���<�y������L�is�Vk��Zaé������J\>�w�c��7�a@���sq��Uq?��0��4��㓁��=����� ��W�$�L�ԉ&�>|6�F<�/�EE�@%��M
y�\���[+�\��ow�8�]�P����j���.7�ˑ��}͢�:C�V�vf%���gq���C�����l��Wϩ� �X�;t!7JoA���Y<�nX�q��8<`��;�p��V]ik���P��#�x�ﳫ��˛�d}rN
A����j`�1-������|�W};�>����}�YBoq����!��:��UT'�<P�Y����~�V{\�Gd���ݯ�E����fc�*��޸	�k�Xg�+i�oR�����p`y�c���"1XB|�[��_���z�H�i<��ݕl@�bЎ��l	٬�.P���<�Ns�q܂.��Ӣ�{�©�s?�3��xiX�i�#�͒�!���^��$:��KU�Q~�{J�dllm1�5����M>ONn�A'I���Ie�M;_��O,n��O�ז,!�u����A��>�+�1�#*��hy����nv\Q�e��W������[*�;��_�Ƌ����#��"���6,=(7&V�7�7�r���%Rl�g���޼��M�K<��Ͳ��t�̿��OftV��գr�NN~��*'��Ja|���K��Y�e A��Zrߡx8Z�=[�\LujD�8���}ge��b(q�ݰ8�:|���/��ڿ/\�~w�>?�?!�U�e�h���!q��M��w����!����>W0����~=����g�j��vLZ�V�2��HԝU�u��ts���t�[�/��1:�\���K�7�&�C�����/������/(�t53M��m'^6��'"��6�� ,:\I�t��-1萶���i�\\�&(�ӊq����b�1<��\kZ�;�K�c�sB:n2���Ž���q�N\��^��m%I ��:����[�3�b�_�v$|C�{$ �@��a���[���?\p�V����8����(�Ǭm��b�N��4�g7$�r�Ͷ��	�s����j�oˉm<�����T�bV����M���ಲ��dG#��TTd�iV��G�,����Z:< ׯ-��1�:��P/?�g�Vͧ�lQ'Do�;�}�sA1A�����>`z��}gx���s��Zo�\�b�AY|>��q��ҏ	�ʶ��t�Q���;�M�#�`�Xc?@e����+��@q�5Uv�-��f�[(��
+?9>S�h�}��caq������2��l�r�!���U�m�n\4����"'o,K�g�η�O��3�q�"y���A���U�O��$��J˒s;[�jȮ�j���ڬhA3��z����b�h�ٗPd ߗ�ἢEP,/���@�3��c{�}f��#��4�)�ۺ��QTჹ؉��H|��e-�*����s����ی�����?\1U�(a�ܪ�麫_���
�YUD�����J�B�;����r�X��U�MD���~�Uo;�D5g�m���t�)z��,y3�U��<y��O�cC��k���g� ��C�A��S���b��n7�4c-�-Q�
�=���ʾXmm@(px��ޙ��lM�̸j^��为�rreӄaSA��v�ڄkh]v���2$@m�PYR{�����' $��r9�r�<fV� "���ƶ�jOI@<u>s	�	��_���wWm3h�ו�SH�o��_i�&<�YQ���o�Z0j��mZ�e��p Z���-b�]ߓ���n�e>��z�[�RSn���� O�;z�L��>+v��=P'��SO~r���������J���v?$|��)X����%i#~��(��M8:�a/�h��*�r[�\5��&�� ��|��G��Z C͵�-�Q�re�����w��i���Oʰ�问 ��|�\Y�׀3�>41��E�tHC����.�ҁ�+��(fIe�᝕��B[NrY����%��Y���B�����6O���Iy�Qq\@
xJ���q9�c��*&Q�x^��6Y�^b}hf��+>�49�rs
dUĵ����}E&�ח��c����FD�`���mm�='�p����w��L��<��t�������Pq/$�4~��8��A�?���K����u+��HU����y�B��7� 8}ɶ}�*�Q{�u,��C�V����ɏ��R�;F{V�� ��~�*~E�p$Y|x�Ϲwb5�F��Ug�]��5~�@=u�0���Ә�1AC��ŧț��Q���1���S]q�+��,�L�%�EI������7��Hߞ���G��8��̪�T�~�eM���<;���r*���TB!J��/����A�7�	͊yܖY�^�����KR�_���  #��ۼ��cvi��苮��[�`c|�����;�|���5�����}}2�M5̓�W�%� �-���͉��m\;�C/a~�T�TPh�����.R[�'$�����m��cq� %�����!��X�3�{$?�FX}��s��j�a �Ϗh7%���9rX9qZYR%�����(��%#�3����Uǣ�H����VӾ}��v�-�b��Hp3�'6�#6�TLq*i�R��}�ں��tT�pk.��ڌa�Q=6����A�\zA���ձ�Y�`G��^s���ƽ�3R���M� �eE;����j�m�>�KՏ�hk:8@��Mo�j3�h�'�/��5��� z.��{1���a�&$���Q�y���W��O���������ٺ��"�Hc�J��>W�z�����lBB�Z��o�3�O��f��/� ſ>��^�D�I�x3 =~��Up�W��q�X��c{Z,?�Y�x6`s�N�	|�"o�yP�[��0�]���wؽ
EY{���t���_׫4=�����Ż����R�)�̩z��x@��K�gz�es���'�I�������D�,qGEk15K�r�Z�.>6O�~?�Y�I�T�����I�y�.H�d�B\��}��y4%s�'X��_z�����RD�HLG�c2}ۑ����h�$:f��@+��d�2"�L��EL��rG��s��$�X�"��Fym6J]9�G�4�r�8���G�q"GM�hk�%Y��"k�qs�|j.�q_����9�h���b�q6M�Q�^�%��Vkkܖ��+߸S�L�~�P�R��1GGV�������%�Z����":��H��W������ �'�֯�㦫U�����Ag@"tG���կ?��*R��`+<��r���*
2:��{��j*t�!S�v�G0jj�-�J�O
lacWH^�N=�����.%L}/��x�ppS}����?x����;�K�啮���Bf�G��٩-�DOiKD����F����ب���i����EEװ��ł��
��3�ڷ�p�V5d�c�z��;GF#v��W#6�U}~c�&�PfpR��7��q- W?�VȮ���J??��(�f�ϔoLS��6�3���fS���ƮR���N�2N��!�;A$>κ��{�v&}�Dq)�8�5xQ��FNZ����lT��D"���	9F\�y���ߠ�Yvt��#B"�ǩ��g3::c���e��PZӳ���.@�E�qW�F���$�L��	��8喧u���3��8�08�8�HI67�֋�p����M���j٧���#���V}%�%�/�*.ɝ�4>��T9.�Kr^H<v���-�o�ѝ&w������b�]���1�۶�7�N��1	'>�a�'!�����*0����>����D�H_/���;n4���qp��:�e3.~���I���c4�H�Ve[���y��h���ɫ}�?�E�|a��:���\,��Ls�h�ũ�	��Da��?4$w�7�@Lc����+{�WD�x��s K�QJuB��fAșW�򡽏pW�Z%ט<W�q�hea�v/�6���n?v�ؔ~-a���w��p1�p@���� ��"W�D?Q�%��WS�@�i��G�u6���?Jim�?�������p��j�r�k��7Mh�pBaҤŗ7���y�ա���"NE��: .ֿS��<�qUd��0�)�Ё�"���CuM�6��/~���N`�2k����5�mcv�&�0��%��Gek�
~���qrS�?%U��*"9�V�sc���:��Ȁ4A ��TӬ7!)h����o�jE,1qTtm���_+p�2�к�U���7���f�?��55��8.ü��䕢ey��+��T��[)��8�(=�Z��V�f0�r�Orݒ���Y�	��xh5��s�y�"u�i���Z4�U�r�����e16Ug��q#b3�H׸?o#?9�(99�������A��$*�27�}��	9�禺�q_g��R��7����s��H��'�m.Me���3A����O�HF6�&.������3zZ��~��fe�H���������~�� ���ll���N���5-g���5@�?6C��-R���r�^��z������A�T��[$�x��Aq����D���/�7��+i��};�$�8H[s}����@W�4�c�@4�߬B.�5��6`��p�����仛g�*��yv��tz�'Y�8"'�zu�x�,���~�l�q�6�u�Ԝlvcv�8���+!+�ጶ�o�@٘W]E4�Vӊ��%��)㒆u>���,��w<i{����x8�-�+�~N�����k�Dp+��U�egB���k$�ʎ�_�P��S�dk��O��T���3�)Ӆ��a4&2۲1��(��=��-��Q]�M
� ��RrQO@��v�F�[\�l��lS���K��tt�Q4�%L � ս��1;D���N�:?�v�n�VR���Ҹ6�FQ-���6�;xɨ�������Ώ�k�O�A$*y˶�kʾ���-f���,���k��.߇�Bje�|`Z5��1��0;(׮;	��
�2S�}/�5E�I2G�jR'�Wyb��N��4>Oi|��ٞ�د������d7W���x �!�o��M⹔����ƸT(�o�_j����RP�
R�
����.���{GP=��j&$L��%�3_��$�	1��\S�~}K2���}�b/l���c� u���t,�t�q�׹.=�l�S�T����&36q�s{K��m`W�ݴ���:�I�+��!��a@��BqzX��e1�Y���B�^�~�`?���L�B9����]�f�f�.vb<O��ST���G>�9+�5V)��+:��?9��&�Ep�G>!hF�v�3�-%�)VG �B/.J_�^��ƈ>Z���_�w$ D���^�����]��e�ɟ6�Sb�ٌ��T&�2Yg*>���1e�;����jW,��p~o4�<u'��{�����髷'�yyL-�Z:gC<��#"��G�鱘c`��
�1F��p�
iBj�-'�Le�,���cN����x����MS���,����橇2�VT\N׮p�?5��K�M2P�7T�-ٖ�re鉘��|��~�.�{�F9I���8�-W5Hܓ�}+m�Z��!��$��u ���>r{^	{�vA@~d<�F�+�DOmU���Օ��dL>=wW �~�"SA)P6���0�����i�A(��%G�S@��вw��s7���Q�������oڣ�Q_��0�~A�z�Ƽq�;�ʎQ���&P>A���R�?ʲ�
I~��w��X`yj ��4������Z����)�Ƕ�<��g2k��zQ 9�9���Λ�GK[;��}.��Q`s�z�M�LUm	�v1z�ӬM�<����0@����[�'�Qj�:��z_s�}Wт��8�*4��Q�3��qAi�^�^�T�\�ǗW����,V���;�����%��\��v�ƛ�6�p�5��,�y���!�N�7n}��cT��m�܉��w<����R�xXE��yc:�ھ쏼�t9�q+����(��	1OӍd��΂�<��0~�V9ⴝ-��߬$F�6T�,��5�;�"�z_Y�����3��pݰy��!�k�Vђ�#h�����x��%�/���1?e3��m����Cʵ�����s��2S�Ҿ��;y����w�>��Vn^
;�!_�>ꍡ�Hb��)��<�:�-T��0�Q'u��e����ըj��vo��Y�a}^$�u��5�?I�s��e��}н@��۲H7��E�Yw�N�:ۖ�s�\����X��o� G(1�"t�8Pr��0���7+�h�R�+�X����������W�J��g�Xw��Y� �V3�l�^ Z�td��Olw�a�\N�6�<��1�(�&���w4�'.N�2��Jȥ%tT|1�0S�o��]��9h�Bl������[C�eeyM�����6٫Qc�W*�*@�LL,d�jS� |����-P��pw���$yluær Y=?g����M�KnȜ�Gv7_�������}I�c�8eC�?r�N����A�G��(�4'_Qvh��F"v"#��]^[V�K#v����O:s�y�Yi $.ϵ"���i�G-���'hɴ+��a�䂪V�k���������o�/NYѳ� ����ul��uR~��́J���9\�^(�XL��	gl�Z���M��s0f(�0��͞�vo�`��]?�v�  �ׯ�&�]q�Bee:��2|�ö�Oh���nq���(;sc��θI�n��D��Y�� �^�HN��J��A9;�V�w�:r�*Qb�´��|��o���X��� �/��E���م�!'��eg���mZ�l<d�Z��C�P��E��j^�z5�|�1�=���D�}d���B7����9YV����?�/��<E��`���̲g�Z!�dZRO��RLȰ�����LG�CN�Efnh��=aGok�cY���='ʝ��u�4 �@�g�m�\�|��� H�01-&�ig�b�����G^8��ݒG���=A�3����Nf'������O��Ε��Y����J�e��U�]�

B�g�4�U| !r]&�J�C�Դx�������()��xډ�x*/p��̂iZ�s�,0T]��Л���ƻ}NC�������j��F)�����w'Hq(���ݵX���C)P���[)��P���{�o�wݿ�f�&�9s�{?ə������c�y�cC�7�@�l_G�Ё��A�j���@�՛W�5ߺ�T�����;@��?q���zfP�����{�|tT��l� �<� ��A�x����n'�~�uv��6	�{{�����[O4��x�D���xy�����|�uP6P5	�w� G�xDt��|y�S�Q��AW?��G�"8��]Ӂ/����$�/|��qe��~z�Z�0wP���X�k޴�M�:	�5]�`P���{5���0�����G����*PUrZ;P�i�p�	�Y9z�}���w���tF�h T���f߇���+�CV,,y���ħm�J�����_�����6o�L���� �5�8�P~�^)�NI���"
"��ԪY��LqX��R,����-qs��N����gX��m҆DRn!{��\���'@�G�>.H7ާ�"nkg��"-.c�9&�Y��L^_|�_n�n2��څf�O"E����<���r�4���=�O`l��{j���*Km�>��|�73���a���	j��B��J/��j�>�.T<>ݰ��Z�~��Ҥ*��ȝ׷1�i�'���6�D�68����x�K�,�;bbrF����e
���Ҷ�>~:Ӆ������=s5꿫kH�x�U�hdZ~?����o�uG�)ӝ�G��^BX��Vt�GG(@� �]�qu����\E������>m���,b�D�9���~��V�X����j�s���9\"��f4F̩�@��\CsG�������[8{Pv� �
�}����n.��P?vG�v?��~Pwy�Dӳw�����o��s�G��i��)�k�=���`v�ųܢ��XǶk4��ˑ�����OPâ�]����.��N�CL$0��ε����'O[�=�������0q��u\���թ�vv3���;��U_$Yɺ)Z��Q��I���&�ր������]�-���$BȜ8+��x�C��d�n��>�i���}��՞3����p�[{f�@֗-s�|�4���!���u����k ��)瘥*#.r8!q<�r��ke���s ���*B��=f�&J�F���� &b/f��ںL���3�1�-&��0�L�|��H������T�:G�p��σ���B�<���z���x����!�vռ�}K��3%��?�T��>\Q�x����B'�&'q���z u�i5/un�oHmDD>!q�J�_�j�;�70�J�5M�����I�	�>k���-�����t,&b4�,e�Pq$�()�(+�pWЕ�� ]�"�=!��X�bgH$�3��b�"�H/�n1��p�j�ؙ/ܚ7�+�'X`���25i,#J���×%0o�/�dJ�.�%f����%�M8H5*ƾ��S�¢�px؝�c.�N#6���N�y73��Bי��5cDp0�~%ع�E� ]̉�jX)��Dna�Ǘ	�ǳ1��^3����ƅG�qn2un�'$��/a�3N\���XF��M"�l�R��ޓwϙ�v�1P�ߒJ����LP7aӎ��۝��[�kơl��_����A�T'$��ډ1q�D�f|x�1.�LcC�����h�=Ž�l�[�ҙ3��q��?H�@LsV���Ưf��@=�&�"�ܶ�� iFl#�����>Ř���G�j\֬��r�`������bB*|8��o�)DD}ˍ�1&�^��hH��N�����+��1�cL�/wT&57jFN�d��0�V��]]��|>�b'қ��b��M�-�9@JMԩ�SK$⊱�	���r���Ȭz��mH��D�������QR�|��Q�0�6@,�<�%�Q-@`ь4����K���VS+d��<M~���PC�Ү�k�߱�ׯ�p��uH=���:������y$�Z�iu���?��<�x�y�&c�G�9�j/~�*޺^9��\<��@~�*,��E'��.�PІ����琧���~��A6�l��.rn�T�RƱN��~==�׫�������UgţY!�h �\�n���4���fl��$����͔V�6��?�4��E��'�":�+WƙI[����/����<�m�PA�_��[oW���q��I@�[1,��UB�t�y$��i=N3{w�p��P�H��t*��ݔށ�.��	zz��v��ν�%8"]�SS}���%1��ؕ3MFҐ�W�o��dz�6��޼�痟i1##����NK���r���)vkn7vmܥ�WU�>��I��ٟGE�����!3�2qk"����ifv4Z�apy��:`y{�,��.~$��Ţ]�UsX'�)oq\�s���9ҟ��8���Pچ��N�aY5*!�5�vt,O�{���mD�=�Y����-�ck5"	h>�d�sOqs�s�bO4aZ�+Q8�4-o�k���I�F���ڴج��!�vUhf�����ccZ��꼺��K$]�����N�m_3��56�3b�����
i@�7�%�$k����̰�.[|im��S�#&��o	ڙX��T�v)���.��׵_;�*�B738���NB�yqgJc�Ai�J��Z|>.hv7�#s �����%�L�����0o+l_�޲�,�>��B��U�q��#���-Ğ+;���t�)R���ˉ[����Ve�f�#�sϰ�NZ����\�`�4E�n�t�tx8q^:���K73^�][���'�,�	̄ڻ
����:!�oc�~��t�/�h���盱�zx�4#������V	e��r�e@��������&U#����5�
�\#+A }��X�x���j��Ô�	8�qc#˳?����@Lws�lt�:��aL����	�YuM��o5��%|f��̼�"�^j("1�cXM��dOۗ���(~��q'-
o������yX=E�U8cpf޺��V+�U��jfRu��a�;S��y�BﴣCO�θ���/�$�4|N�&F���3���[K
��H�����%��G~?��z��GG^�{X�Z Z�STn���,g�$
L��8�ֿۑJp�#~��xэ�%S泋)�آ�>f�D�d|���60a�&�չM�񨒻t������?�muӱ��p�m���&>LR^gmHO����N:e��R������B/w�������Ո��_�gz��S��:t�U���ß�y�Y����><�u�H�ϱ��;���5�J�}-i�#%���
CC�%@0�]~n�.y*�UA�bP����Va���P<���Z�kp[��������[!^u�� �+�m��팤^�V��#�w	�y~��a��y0���ZV�G��=�������;�3 ����j~'v��s�%H�}Ɯ��6)dIr1 ��ϟe�Y����q��g-�lx��l�����8un%p�&�����bq>(��hX;�M�t�ט��ak������~܈a9@r� � y7Dmh��e�|�C{;,�E�s�17�r6�rUl��QF�߫mh�l�t:D(�*�4FFSY��|�ʃ{�^k�l5Mf���7�ɶ�����* ȑd�Q2�"���gY� �e�3�>�R��?���0Q5r�~��?^ړf�V��^��I`3���8�N�d'�)�n����ME�F/�ᬊJ�
}��l>�c�*��ȿ%�T�Qq��2�DƮ�U�x4X��������a�|�D�yr�O�I�J`3��:�K֞D��/z��W�b�;��C����C_o�k�����%����'F����ws�����
�K@%_S~�C���a�~m�$�����<[��$�S���k 5�-И��TA7,��^�� ��4eC'/��sB��e��ڽ�^&Z7M��mss��,��w�ڃ��2ܻu��}5Z?,,�$��]�C�,+�D�Ǐ���j�ᅤ��e)�ZpjMV����yM'���K��\G�����e����i1Me���A��)<?އ�w�Ũ,�$���^ҿX��>)������rh�!�����=�=�=y�>+'b���7pQ����p���tf�%A���۟��H?�ȃwvn�1[� ~��h�?���D��]&5���ш���,A���h��Yi���z��t��+�Q~�i@ď�˷p�/9�t퉞����\�p3U[*��_�Q��k >����Ma�R��t��G!��˭$�rz"d��?E�o��W+��& C���X>OO�ey�m��������w?_o�����u�a�k�� j��Z�J�H�[\�1 8b����>U�bɏI�@: X]�x���9]}�"
=E>|g�m�i��W�(�ׇ�?��8@�����4\�P���玽��������k�VZlֽd
���הOz6���z�ޝ.4�,B-��H& {R�)p��l<dC``�i52�d�[��^����#�xÖ�Ҭ3~0���գO�x~�{C������;e���ǳR�\H�4��A��7�b��#&f�o_�TL�F1r�l>B3���18���.�3��G�*K���W <bI��)@,�T��b��C2˽Gš��q�k���PM�m��	��HU�"�����S��V4�>9����浯�]\x�'����n#��=�m�|�)ׅ��ހ���++��܈���ڳ�l��6�s�c-5��Ƭ/;KR�	�� �J1���~"r���٬Nu�ֻl�y����L<.�/����{v(֏�;����\��_n�b����t�6ԩZ�<�g�?x�����?����֬��S��Ƈ�
���S���O��� �t-���B�zW���5ed��N�p���k����{�"O! ��$	����p������z|�FC��c�	� e�3�p��L[D��h���q��,��b{$k����<�j<_ȯ�L�����c��e�S����K�M�R���Q῁���}Jgm?���Z�ލ{�ț���VD�x�~]a;o����E�՛��е�8�$(���k!@Xәdht�n���7;?2W�Ol�Ǉ(��C%�ɿ9f9�j�Ӳr��6>۰0�9� ��z�%	]��ҾA��<j�݁���lqW�`�ӱ�8�A=ּ%��f���aƜ�Us(Kh9Z��|obc��η��a���OI�	�k��3c�i�1U��P���w�6��)��)�й�QP���|4����\r����M�Ni�Eab\�gR�`�1�%Λ;�S+�հ�f2�.�@�p��͹�:|9�"W�6z\��kR/��pC��q �}�b��L������΄]Ƙ�bP�$��/�?�A�4�iKl*?剅ŀ��כ?��a�'���S��LT�W�[�7n�,r�DF�]����} Z��g	�2��<.�x���57Ԗl< ����%X�� �}	�O���~ =z�h�Bܤ<:���ŀJ��=vQh;@�kO�B�k�Z����Kf�[[[c����P10̜�1�8=Aޅ�WJ��� {�d��)������UZZzuS?�] -a 4/�
�
����{,��ib��Cqwlf�AT�V�^#O5������T�l�M����"rd�{~��a��"ɦ}��ԙޡO5�2k�~xxXUO/���?G)I������4ln$�`��1��.^��n��)%z���|MM�+,���\�A��&$'����LQ��]$50�K����Kâ�����Q23I#"'���
�?�S�k��3�@Sb�a��e�]�Co;;�b��@M��%t<Yd��fcL���������)��4m��|S���<Uĕ�BB����H��C�*��[a�p�!�Ï{Y�_�����eh�4�<bOG!�߷�԰���Bqp����� �_�L��E�?���fՄ�KK#�>WS��SEK���i�曷"��2JJh


��:��ﮮ� ܘ���7<b/�)�Y?Yv�%��?������������B�(gu����M�P-�"ɏ����"����wn	�X@��E6ONS�¦�T�p6gW�W����Y����H��[�յ2���߱?�Uݕ6O�[H�㟾ڔj0���3���381��e1eͫNTka� ��Ķ��@���O!���5txX��Ç��:\b�ۢ��<�����D�Q{�7$h@Nى��͇���:̩ȟ?�i��?�L��U(
Yqh����`޸��vi><M���� ��v�]|�TT�b��P2�/V��L Oq	
Z[I�B��*���c����Jڬ-<�hk�\K<z$���Χ�˼�$-Tx�,e\||jBTjl*Q�~ǹ�#�])��E;���r�r��ml ���-k���;�p@N���i��w'�ryF�Hѩ�d�4�
jj��RRRZ���eޕk��?��Ph��(ſ3�W�����ө��#EGpRZ�%F*̸ZgݣŻ�D��]/ �w�r ��e,�K�oJ�|6F����v���0�$�HM��B�
f�RQ�	��Z��U?��'�EE�j�\\\L(e�<�7p?p���:j��ӧX���0�����<U�_�]м�ߏ5�z��	�kφs��5����ƾ˓&�?��π��i`�I����������-�j�Kf�8��e���C�o;T(�S�R�K�C1�j�|�4���˗��������@�X����hyZ����@���_yu�"Y;;���M������KU�t���>@v^�pe������z�����U���6����@�/ұ��5uM���bzSH�%`���jPw���&��<U��%��{
��e�w�_舉�U��ER�j�9	9ED�y�>�u��� F�Xq���ݶ\��&9�+�;z�0_�,���KL2m��&tsq?c�c�~`9��^QG8�ڇ��I9*����Z,@�ׯ}�-g��]����Y���?<*K�Hn�yy�C�*�'�A�S
�Ţ�OϦ��7�fB��	o�:���}IE��֬�0�W�9e[�����fV�/��TY�f���MF���^���,������U4	:e�Ɋ�⚚��[W�d�rE���a[�E�SE�/q��1.L ;+>JLL�����:�2�\�{9�!:�ew���Y �tj-��<ŬPz8YYæ�i xu��/��A��1$��,
>k�t�"�"���2 �rEjR�����o���d�;֖]\WiK�і[h��	><���&ʙ��/R�+	.��)��2>Y��4�����O�-=K{����HJ�)���_�|�Xc��KNT�6�hc�T9�L 2M�K�zqMMT�B}Xc�S�slo�*�-�*������K"��.�2�����F'�Hpc�K���Vu`���Y�2ޜ���C����+͟���ڛ�����\��@i !65�:��	 ��V�S�W<>US��3�fr9�7���ᴶ�sp�X����֧�h��΢rtqS5�������kU`K�2��t��xOr��~�݆��JY�H;�2�G��5���|�ɑ��:���Z�	]�������4��qY��Ī�5z��"��Γ���T�l��vF�~�-��|�a���nm��9(j]��B�B����j�ЎU��;zh1.�_SSS\o�&�80)��?��#��C{����@��P�$�Ic�������Gh	����ɮ���pz�e-����2`�-�49��X�r�Le�j��kd��6�:T��:&T����1Z# ��
���t{�٩1/Q�V��� O�j��[�Wв>�S~�C2*�ƣx����1Z��h��;�S�������k�c{���a�n/4e�k���%(<%7�uxWU`(w9��<�# 0�Hjͥz{g.DG=��#��̙)0��n`��MO��s�����}�V���Q���2�| #��,��z��dh0�`�3P�a�*��l�R*��z�AH�ż�p�-q`�B}�!�|�)>���zF&*�߮�;�_q�Q����G�9,����T�'��yM��D�,U�yo�W�W���$V2c�3�*�_@���Ӏ�=&�ɸ��ڏ����3@��n�-Y:Z��41�}�m�r-]P

���f^s����&�8F��J�yfA?Ө>P{,�X$Oq�KYl��Z�4��ۙ��b��ZV}V�ID�e5r_?��]�nmw-Jձ,��[;cƝ��$Z:��=ǘ�\�{:�C�����S�T�7\�F'��_� k%��X�%sک���4%�>��)dI)c0ZId�q
]-������߿{i�����H��G��r)��w����by���=�[2�j��R�S,�2}��[�[��Ǐ(z�F�OMr���ɭ��Ť�%��_)���%��h��Xp!�ŉ���rd���˽	���@&�{b�P��#	���47PO�Gj��_8ɪJ�$��zU�"6����B�79�fh�\��;�����@Jt#&!&���aխ	��H�')������ef�Yi(|����y���+��{Ш&��^q�Pȓ�A���\J�Zyii�����S��(m�'ː\��>�]U3Bx�4�$���@�1h���ph/<��wG���[oT��eff��S/#�i�a�U���[9	��<�{�ʒ�Z�8�x����t"��>������H�i`��22M�W*�M���/E��5:�����{��Y_��* �?(r�m���̟,�P)�գ&�ji����q
RN�%�,�h�.jՏ<���3�G|@3�=*a3���l,p�xO�u�u�{��t>5���Ȉ�B�q"�B�>ӊ���5�魄<_�_��m4��^�ڢ�܊�#n��'22r��na� Զ}�9wޏ1����@�g~(�%���Q97oM?��~�P���{�`,>[r] �u����PZ�T�z��Uiu���/w�h�������G��]�w��c35TV}���!Ȅe���@�R�roӻ�`<���������tbA���f�h�@a[��'Cv}��5~�Z�����9,�J��)�c��(U�3��˜:��sGp��!I�fC[�A�?�����!��.��z�Sr�)�	(n�O���^t}���fJ�����'�I� �;��&3�!��/��m���	7�v<ǉR >�Ѓ�S�E��ga��h�]�
�\�^3G5�!�9���5s6q2tI{@���
���Dŋ�b���G�-N֌K�NYG���B6jt4�N#��c��͚+���7�����-�w��T�^~Eii��`1�E�Ħ-�|���R9��KV}�p�^��)-������`��ܢ��̨���=�ki��}rJWƘT]���b�7�V _�V�ɿ4��T�q�����WU������[�ރ�.v>2�n'�_��� 	\��!!�mY�������壖=����j���)C�ܼ�8/��+u����|�)R��&���y�/3��k愹�> �q�p�������5F�`��@m�r󈕮W�7��3H�K���ۃ�w�h^
�~�^�%�"�M���&yQ�u.��U_�����|�L���	��qe�������Ǯ��ؘ�(w:|�,�oOǲE���#e?X]\��f��g��f;x�{��ms����.F������<}P�t�@x!�#[�*�5argh&gD���v����-X0�)�
� �N)������U��V[�wZ���xو e�	ֹ�B���O���5�BQ��/3?F��s���I�BK�������t�
4P��~Ys���8N�8�1�*�Z�І�Ҟ�F�r���l!Vm(���x����%����Z���D��>�_MU�_�m�kZV!ᶐ�B�J�U����|j���d�ęD�N�P��	!
PF����֢�ܓ~4DRI$��T����|+nK]ڨ����v$�ÉZ���Ù\K��d����i��^�{ߡ���?��l)�����}��-�Rc�?b�����[��\��v�'���9�n��=�O��6q\pb���]ΏBA��&�N�t:2��:����Ȕ��H�$�͈[��7ԩCD�Y-����vg�i�L�em���1�qY��K��&�%+���� ��Z$��Fk�۪�Zg��{{���9�=c.��n�"5ϴ��4�BK��G���_
o�WE'�������e�=NX�*�@�宕,�p]e�d+��M����/C���k��H�EB+Ф8��ټ	MyɃ����н4�A�S����Ƣaa]�{ey)���0hqTp��ҌG��'S)����WQ��2԰jO��=,;I	>�۹Z|�R^�u90�RP8�R�B~h��d�u͌0b㏥�����D�B��^�49Lb�K���6Rd:�{D��}¹�j�ҿ�/w�K2��¦��C:�uE�$r�x���1���C�S\{���m�����-��󹉖-#O<kA����Q�6�#�L8��]s�`�����R=�x�ߌ|/�6��M��݆�~�|(�9��zjU�ܲxf�]�a�x��c.G���H��S�6t�/sz���C{��٫@���7�O�U�-��R'��M�J��?��?��`�֐��>�%�"h:�j��"N�V̀�4<��rzn����fŪ���i	���
Wbq;W���w❄�M
rd���Za���-�_�3WR�g��w�e�O�fP>�c��������!T��v$�M��f9@�����_�\X�HB�Fj�$���[OSj�x�!&$*�d9Zs�_}�\�U��͈Ѝ��1�����W� c�*@k��8z��(�S��B�R�~ػ�2^��ge�"�
x���b�xzr}u�Z��ɑ
9<JH(����{������P�@���v>泌��}���3�o	X.��Ɣ�N�5S�1d7�����79	��'
��R�"�����⸠�������8��c#�)��:3�f::ƿ�d	�S�m�����\���/�Ze E�ȹ�}S����!��u�f`������}�����ަ-���!O���j֟fnCW;�o|�j3T�a��Мg�6��딌�yb��i
-ɥpǞG?t��z{�.5�4+kJX�Wy|AK��/3�-�Pϲx�9���1F�«�{L��PsF�:�b��<}��*&)�׿�pP00�7D��5x���;�Z�a�-+�@j�7�����3s�_{M�=��M���-Z8�Bw�XAa�������p:wr�h�L���0�.��p��p?�x��2����r���3������Վ��������ǃ<PÚ��./����E�*��I���/��D�.����_/]- x'�y�?ng/[Pb�35[z� �N�8,󖕐8&�(�BPW�8`$/�)tY�UP�*�ے\ZV2�Zqp��>�����,t�byW&:?S�Ѕc��~�'B�Cw �	�Pc�����&�6H�(q
�Y�@A�#l!� Bs:���;�r~�y7D]�W��-��� �H[�.f`0}�>�2�6���p�h�T��a��P�F ��4E�O�k9�ټH����t)��r�(ZJ�/���'3�#�r̹cp�Pes�-$P�4'i�	6q�Jb!����雜v��!��jԷQ��^|.�EʰX	n�ƺ���ϙ"�r�|X6�������IrM{)���.�݅�PM�1�чmO퍌(��V�������[><< U���"t���P�n�� 	���*O�(i�
:*����������]9g�Q�{��R�h"�"���Jf�6LP�lQ�x�@���o�SfxnII�U�f^�B��>%̓J���v����l�=1z5e�B3����T0��Õ�rQl�˿B^2w��"""���@&d"�O Cq&��+�w������Te\(22U0��F؛[j�;�,����P���| ���{?LY����L�G۫ʊ���e`+�
��>y�(�r2����� s�o���d'��h�&���L��Ժx�NOw��(�[����¢�4�B����+����e��������bK��Mʩ���-O_��Ǌ�.�Ы�M����������tvvm+�

DE5��5/�e��{x(�����a�����	&���6t��տe
Cy�~�ƚ|qyY���J�?xї;�։�*�fH��
����X1q��q�t�,k\m,̒�����}�sO�e;@;���8�:��,Е5M ��sQ�g�I�����9��e��P���z�2(�qru=?ߛs���n�ɣ��bz�TL��Y"�%,]c?B.�UT0����x��5[M�ra��̄��5�[�D�l�fQ��P�`y��JTzs�1�e�(�=п���2U9m|3�Pl�{ �b��o��'z�(�p�JC��{���g �!�a�dP��xZ��.7z�q�����-�M��}�[�<>�K���3J��D��'o�OH�N�9�C��������ዴm�a���̪�r�	W�L?��Y\t!P�Mo�$�	����/4LĪF���+���WW�i3_��$���~�Ǒ��H�/R����ʷ����9K�`�=wFePNl���s���0�`{{��A9~�M%�vF���Pc�t��l(��I�K���Je�.�9^a9AC�$1���KY��vk�PR�q�N������&y�p���k{"1pt/������yɒ}�����=������pP^ľ7���h���ooqH����wH��ԏ�.�-�x��QQ~%��+|{iz�,��9ٶJ��7���ޅ�l��gj*8��ڳ*]�@���0j����cz��$e 	4��6��Jz�'�D^=>[;8���~��O�����};��.2���g��uN����PR�VrE����0��аd���1������ZTt���C�yRwċF^�COO����Z�=e�j1IJLJ������q���C���O[�k��$C@'��&IP�v��7z�βA������E���0%�m�N0eG���1������-��	�&���_����X��OM����42)�~�<K�s?99!$&�~�K��c��⩂͂��������L_-^Lķ/��ñ��;&�N�R�$��A��خ�(��l��o @:��.^^)��~:B22����%�^�\
�}+v�X��la����VV���HE�O)���k,B�W0��XC+::(��ؤ�.�z�;��- gED��	�?�Yg���^T�+[�pBG}	���a�>��������c&O0[k��e���EL��mک�_�la-Z�ͧ��x�!An�WJ�d]���;�<�mZ�LJHHYi��e&҃�Z�
�	:::����d�9�e��)3@{�H0�������PK���;8�̩ݓ���./M8	�ڬ@�36u��74�ߵd�V���*NQ�j/UR�2=���&$!�:tf����4 7=u"#ͼ^�EHmYQh�m~�Cd����T����	#�[,n���e'���KD��X�	�y?��ޗW��]5�222�Z�I9*�Ol΄���t���+G}�g��//� Ǻs5l_YnH/�h{ɕ��o�O�.����_�G806z��i�����K��X\UF2>�x����~�ymUѲJY��m��������9�T^����g�Wf��/���bũm#������N@V�%�JSc����s)1�D���d�e0D%�]>>Ϸ���$/D�
h)�}�5����3��1�ʞ���yF��/D-��U�:\�A���U���G�䬍E bb���>/7�������)"���wDq�.I��l�-�[�r� �'��	y
,��_�C��� �G"z��9���/�cvUh8�� ��ܞ��7R�"���u��K\1�M�3Dz�.�"n�K�)gz��O�a	-a &c>^F����?��羏��b%z�s�˯fO7Y.�b�Uj-��]�dfpb"R�+P��c�3��k��1Y���h�v/Ѡ90"]_�]=��*ggL�6r|�G!�����b	�/l�]�L�x@ 6���F���s@\\%�@֗��qZAѦ�����V����19�(�f�Lx�G� ���_K'!�2=�"w�0��nP��z_e?}�u��M��w��#Jx����|���-�]oMH&ش�fxx0O��`� v������ʕ����W,�(��A@o�� �2�Ҟ��Rc]��Ҥ*Pqp$��ۺ�bGbP�����jqf�ah@:E���9����+���ޭckkD�,����Ǡ����# �r�y�R63#7p�(,a�,���SE�R�.���ո⸽�#^>�� u�'��@�Z���s�5�&��g�	Ċ��v	�89��yc���S��������B�����J.�V�w�HO�jL@낤�A$��/�������ʘ��>��o+��_�^�=�e��/���g�.X9ykZ�Ҥ�_�*<��������/_�W�Fk'n�Z�p!�C�=�����M���/6y� �L����d�|��FP�!OT=5�B�8��A8XR�$ H������{�/���W�x��bɽb%��t9�u�&N�
-�c��>����n���p�փ0�Z�ǋ5�;k:f�����|5�s'�B�̩�Ȯ�ՉT�o �C�u��c�l8#��l�
�\���pʊ�gJ�F�H+*�	'o����k����DKcʘE=�{��wb�$$%��oo�T2:��[��ʾ��7D���N�!k|~O���"""谐�e`j���6���g����pzB�x�Zn^���)�؎�`j06m��.{ǳ��;Or�h�M aeO��X�t�: �Glw(����p�@�� ê�RvR��o	Ԏ��J���>K�BB��K���t��@2M�}
'!*[��/�X���u��][o��Inu�_`PC���NO���8i���!m�c��Y�R=e�j���F���}����?��u�n�6�){Ŭ������Ъ�b}*Θ�@���j1Q���V������@ԉ��pL�ޙnl��|���O!�����=i[�e�W/Q� �'�6뵻������l{�m�ed���Kn����r�b`�<^��9�-�4��733����]*5f���î�83�3��-�����Xک�0B��)j%��VGպU����G�H�����fq�Y`��a"�c���zã�	sv���C��~ڭ�D�Je�����y-�GpX������
$ɁF{{a�r������V�i��O\:gEK�� W8�"��@�#@B������>�-�n�o@�n��T�y��Gb0�m=1p1�HoooN��=��jRtL��3SS�_X�#�I����s����|�D.!j�sƜ���������5�0	*���gj2G9�L��0kv���O� �֞(�y�������G[na��X�b��{�P����҃;[JNF�+[OM�g����0��A.��R�;]�z=ғ�<)�Xʾ�Q�OY������_�_4�ݓ��kI+�[�HMi̜*��bŗRn/���ڔ) �'L�dV@� ��j���9`�"Wf�o`�$0=V����ɠ��k���8,T��ic�Ծ�l�
p���fI���xdz���@�>� ��#L�n�΂v ��Ƅ�Y����
E���
oiוy�P���T���?٦�*���R��yW
������⌘0�~\5�a��{�V�z��1�}������A���%3 ��:����ox�>�%#M��ҧ ��?�:�`�ֈK�8���b�m]�_�� F�I���KVh_��Tμ����b������e!o n�B����9���'&6��T ����_K�jB��0��R���h��'�Eʿ9����7����T�E�[��T�͊��jpT���|�mr3,/�����$/=r�'/t�j5nCD�b���'$:�A=�ɚ�g��@E��D�@����j�/�[�Q嫽/a;Ј�K�|����"q�W�.�9+��>h}�A�M�5䴫}�샾�o^��~�5�	�˒~�ՙ���wS	>���Աs���Ǩ���U(ow5ھ2�Wʑ}���v�
?_�����,�b�n��엻j����j9����l��������nX�H_�J��d��\������(J߽�n�9l}8D\�Mxbd�/v9� <�[�r�����,��_62�

\hS~�*���,eu�v��⠵��
�����r�B���`�u
<��[ᘗNŸ�L,,l���O��Q�O2~��|��$�j�	Z��q��6��g	��-��Q���4y��o��Ǘ�J��dy����l����$G����`�w�c8��{?P�&"�h���79ϭ��5�V�x!��3j���L�c*[l�*���N�\=��"?��B�'��.N[���\�,�i#66�V���}�辎	N�'s������|��F��Xͪ;v%bqr��m*i�2����н�#�|*���`B#9η3�>��^���緖��k�:a�h�T���U���}f00&��/�[��G�=�#ܦ��8���[��&�[�^�~���{B�Wo�"*���ѯ��{���;(������f��İPtsXw;���HK��์�PS�0�̉���ѐz;�4;���ԯ��!^BH�G�d���A�%� �(S7)��DC}|������5�T`[ Ȣ"�}v�ր�Ǻ�� J���ɘ�Z�_�OW�V��S��^)�v�V��X��%e����*c�IԾ-�SaA���T,���0DK,E�i�j���/��|7缓��{ν��{�������	�N����2�0�в\`{�S�k;�XO�PHV����CU_Yx���]�7j�a`��N����>[�8X��;���eI�3h�n�AIF=�N������)�ݕ��r(���(Rӆ6���*>B�,)A�;��_`(�z��R[�t���&��9cX�H�l�yi��I��!�V�l&�����_����=2u�KTW@��܎-�T�qDi	Tv��V7���3X&X�s�j��{���T0��Ô���S���)��&�O�s����"�/�5��?�	��P�.�1��:X8�r�`�e��_��ηJ���g!��S>5�UUr�r�T�m�mv����"�`��L�NNn��Q�y݃�����j���gCN�d;�~�#9�u�sUE%:�������Ǖ��Jg��d�s���j�p��_����Y��O��:����S�����xa�g|�{X~�ϕ.�������<v�[)���3�������z1%.�0�2��	�yТ�tȣ�V���}��K%/���>i��!)������ּehB1�(F�Nx�e�PYy�F�p�SF�V��p���"������xk��.luN��k:]ؾ�ɐ�u����J *q�Eܶ-��F�y���~��<,)&����4B������E��B=)q�.��Qa���Ȝ8j�<�4Z&z���4N�[u�@�����1��?1;^4��֮�8W��n�19�\��Х�/E�-y�e6���=^��9(dbG�3n��� ��б*IV��c�J ��������2 v�2k}b���������H)�̯�i�4�Q�m	Bz;����T�f�U�,�A��k	H?>��AUM����s�&�G��|��i���?:ǳ�@)�a��l��������W�Z�z� ����O���t?��̚�N%��KtV�����lr*@;U/�G_?4d:�|՘���+�����Lؿ|���b�`����cu�u޲r�k��ֽ�3H��3-��_��e�%�����f�V�+8m��iU�D�1:y����_�Ľ�����VƔ�vj!@�LS<���j�+d�DT�����"��
�\��B
-n�AqK�d &�xSs�fzX�Uk$�_�x�p;}F�H=���"^'�@���k{�jz#���7�SM�qnt�]\���Rh��N�E�kx}Y.	@�Y�mo?��0���ؑ���WLR]o	��~�n%~KD+*NMD���f�Z,q���IP�	0������^)E����E��b��𵐒����5�o�I{��5��!��xr��܄">ᘸ\�ksd����b�sZ2:��c!�B/\r;�󝳞��͵~��.OXgr-�O��ib*�V2�c���Xڤ4e�C����Q���־�����^��$.�1�o�qGa��O�|�?�8RC��}ڈc�j׭���l��}�����O3;��	]I��|��ܫ�\�h8��t���2(�T�WBO9ak��&��-ش�S�N=/���Ib'0Jp�^�˷N\�������Q�����I�Da�ⴥ�#����4Cw��\�(�y��QE����\a`�cV��#�2����Z� x���+�@�n�Cn��k�M[��X�'d��Tx��{ֺ����ϴ��q�<~$
v�/8��Rj'����џ��D~JRqR��ade=�7>����������nc٦w�f��*����Oݞ_
���5Rۮ�W!P>)�Sp�g.r�=� �0m�An�_fm�Qv3y�do�v�ָ
�%|�]I^��Л�{�u�OSI��ӏ!�
/E�H�� �r�:���*���B|�?�z0�Kh��S*��W�z�?���q> �(�ٺT3���|���a W@(� �\�����+���z!n��Ъ�Ppd�m��$uX�z�3d���ù�A~�D�kX�
�^��ݗ���j�},��C5�}P�ӡ]߹�@�{cs�_.'�Hݲ���G���h�U�J�V�q�Y�s����F�
v�m�d)����i���A��w=�0�����>Âϭ#|G={��;L��v�<�]��l��orVs��6? =�7��d?lʲ��"6_W�e�'�f	��)���Y�m�{pZ�1Ҭ!�Oƾ�p6��6K�G�ܖly,�(LMv�(L`w}o`�W�w�����~S��4m���kcʢ���op%���l�����ϥ�Ln��j���R��(P�T~	_����P,R�����b��a�g+�7�⍉�&@W	d�V|��oځ�	�] /G>�搈�mUUѣ
���������qp�i�V3��"@���/k�N��96�1�t�<w�#>�o��dg�C���}�:@�m;�����B�"E��l��H(P�����P�K޿j
�w�tBF�]F�9�>��|���ڪ�TB�hR�:촌Hz�����	�s��8@�(	P�Mc�pV�<;�0R;o���Yg�r����%7u�W�J��׮H�B�"4�|)4��bB1�OAMF�>ٰ&M��^�tγ���S�ã�̽�e	ƾ���~#��S��y���l�5��v-H���[A�2i+<�@��a�4e��r0�B\	Ŭ��S�^�Y��&&��|d������q���O4�&��4���<���F�.wL���E%I�����=3�3�g�2/��2�/�6T�[-[1)��Ms-�U�x؊ʤz"����獵��X~#��en��Kh�����<#D�⽵})���c�Ũ_�*Mfjz?�:>]��pq�?٣�B��o�L�C���4�Q�P�����{����:�kfu�wN����ݲ�T���PK   Th�Y����  (  /   images/c33d050f-98d7-424b-970e-349228d04709.png�wgPSQ�-E:�BG:���`� %��4C���!�@蠡7�(�B�7�&"
H��p�?�{g����;3�������k��白�ƆnRsR����4%""�Z%)!�b@�1�\� ����U͸9yZ�?�yJ��@w�u�!�X��z@$�xm{`�7������w~��69�����^$7,���[$�靍��D�cV���5�Ь޶Ě��07�8���49ehz��x��=�O����*���>��jw4�l�\���G�|�qL�L�B@�{w�]"��/F;���F~��5FQT� 
�������r��M��{6 ��$56>'NQ����5�.�(\�uCb�+�Y:I��#sٟ*�l��sڇ�5�����:>-��;[i��=6���d�cO���R{{EU ��A78j���#x�Po���E�h�t$m^1"��[�9���z�����������'(>s�nL,���ˣcg�֌̛�Pܴ�s�ovy�M�z���g�}�֯#۴J�;wf_�;yDdƺ<Ԇ�F9!b��x��.%c��X�0C��w���ȹ#���xT~:�����5�<q:."".]M5�Т��4�E��rҺ�d�h�g��nU.Q�	��Cy8�y�ef���9ɖ�7�Zb������=ߥ�l
�\���e��y��j<���J�SIM?c�c@CD�lb�)BW[�.�<�_��4�f���A9��?6??��i��vS|���N��K�{�Mb��U�����=l�ڃ��/�"8�s�����h�f`Zضk-$��|X58W�%�����ɻI�X��}U����vW����3��%Su���w�x|�`d�F�z�ߓjӍD�̾���0?�uI��d�&�DQ�D�M$����m�`�����ϭ��'xs�LP�/G�-�vTOT�Yp��e[y�6e2���Z��HE�Q~�×������W*�{�8McxD1��U��_}�A��U�ɟ0׋ڕ�bS"rT�f� ���ju�#=;�ذ�IO�w�Q��8"�Y+ʅ��2k�[�K%/�	HO�����v^����dv���j���)�F��:Igax�&iD���ܜӭjfU�[�8�.�]�iv��R'���s�i�y�a]q�����M�r5`_��Z���jg��pP��y�c�y`�
}Pe\�?[0҉lyT�m�ow�:hx����(��)�bÙF��*������Kh�k3��ƅs��)Q��4Yb�`�w�]��4���~���Gl9�c���.�=Ɨ�O����\N1�N.�{�SMrM�M��":���i^��p�࿉�Lۦ^��m]RG�[6��"�i��$�%��)� ���>�~2�S�w�]���v������l���5J�4��&4�n)�IU�b�s)t��r(�c�����.�� XE=K+d������W��bo���Z�M_�ܜ(bU/$�"��g/K.C���An�3�n���o�0�&q����Q��ݻɂb�;���C�4��@�ȝ]Ś1I������z�O��ɳ3�p7���i���b�����f���_?Wr�7�Rj��^4���]<�T�yj�{�g�x��G�����������������Q�G5V��P<����3$u��m��=��{�� vm�	���,�{$�S�.���ED���f���ؗ`X,���^-X	nث*�r�~��`��/%��{�]�ץoߦC�펷��g�����{�dƵQ�Y���5����P'���+��+���:�������֨m�`�5uo���e`�<4^�����r����^��g�}�ėM��}�c�Lb'�_��ޅ(��n�HD8C�O>�-1�beS�m���?}ߍs]���!����-�f[G-�%�;�s��2��pG�7���%qI��w�2W�u�<��1N�Fhۊ�&��o1�f)۫��ٹ����
����W��;��Tf"�lm1�Hc�S�Y�Z����0/�G�C_}��f�g{x_vH#��/w����l �q`@IB�m������K�G����?Ɉ��X�t���3ʯ��H�*��4��; 9/j7F�,����!A���<ON�����-Ӕ��c6D0]�2m�(�ɘ#:��^�Xk�|��JU��⇹�;�x!�͜�����~�"�������$�]-��|��W��T���̪i�l��_]�3!�x+Ǔ�/=_Qm��Y�ѭnr$7ˎ�8�5��h�}�A��~�sw�ֽ<�b���*���7Qb�&<�DOA��;3�T��H3nͽz��酓�Q�Kw$<�HQ���І�!MjM�%'p��ʶZP�䶗04M��E���QDv�MOY\8��W���<�����h���B]�T\��s|���V}e���
o-��^f��#Y�L���[�ՠ�)��� �!�8�u`��#Ϯ�(/�L3�~c���l6h*����� ��xi4|YZ=��.����I��**��ȜXC�n=4���l������m���Z�9E?�WV����g�ۏ�+n5�i�?�ZM����tgB7}�ݕU��ǰ�@`�R��C��6Bj���4�\��.�����z����}�d;;�w���z)\����i�}rl��c��t50ȯ+Z9K������6b�;Z�=�n�R�^b|y��6�t�ȭUmǻ�#b�˩f����̿�Y�X���Rh��Z
@�A��!�0��.�O��777Ƿ��ԫD�E?(��uPs�4n~Z\�9�+ٺ���3`�2]~�W>]�.��gw����� �E�Ҟ����QL����ڝZLD�y�k�ȴ�/���������kL�/uA}��^���u<E]A����
�}�G��PY�����r>E�q��\�/^!��?M��-ݛ�c���V:L�t��O�rbT�X��a����U�Aj`�U�>���R�J���p����ߣ�<h�����𒶫(��r����+����}F����u3^aI���L�S��q��e�F��}��V�q���D�(�9%]17����x0���Su�#����_���@hg�oُ�-K���j��c�QL�����#"��*�퍩 }�OO��+�zl=oH��'���_��/��`�=Sj���e�j�_�ˌ��^�r.�`���\�����3�29�����J�=��W��q�#ҿ>��k��3��r��Y¿6?�� ���[��ՙ\(X���d/��R��\�`�CT@���x��������n�o�;Ƚ����"ǝ��z���ܛ�Vf,O�.���F�`���o9Nk{'1�����S�ǓRz�dn"�2�ԋ�JX�"?���qNQ�NvhRG�׽�%A�ѫ�h�h{���J���8��e�����|8%�hܡ!�^Q��!����|X�ť}�	K�h:�q�٨0:~dWg?#Y����(�E�YQD){N2������ �3?�p2��;�h���o=��M�v����1�n�n}d���G͒M����/�Aۥ"rW�$w�yM�yF�>N7�Dm�<CR��d�A�E��0W�l�\��Q�onK����,y �g�E��5�֖�U��a�]P�M����M%.X7|=j��E"Xz�c�c `�m���Ͼ�$GL)��W�w	6�R��S�
����1h��h�Uj��#�/o~��5d�����HN&�1zJ~m�k'q��װ~�  ��g�}a�g�V�1�pͦ������%?��%c���7��u6ׯ�ܼ�,��L�M��H���mI�4m?	�8���a�QSф��b�p�;�r���$�'��D�S��2 9��Ҫh���]�_b����;�U�E��a���?��m�����?ͨ�6�r1����Y��  ,�}W��X
n��u	�5��(�C��*4�t����<�
/|[0ߗ8��@x^px��Ko�ŷ��}) u�ܽUG����&����9��#X'�Yrk�1�􋤡U�0�P��;+VH�j�����}�)i���!J�0�B�¡9��7u�'��P�t!�l�n+ ���K���ؤ�0�)����9���'�|dE/�Xؐ�/Ґ�W���߸����:+��#�:Hs?d?�Up���W�*3
����1���Ի�XQ	�swS��9y�n�>y�.Fp�����5���k?4�����?a:L��!_5�;�%��t�$������&1��N�0�
���~�����^�j5སZ�P�QѺ �^�K����}�3Y��@nw{l�,�!ſG�5/��5�ʛ1ͽ%k]��ُ�&���%ߠ�$�7d��CU��~ע��(]����q,�k�1;���^���YxT���<�#�v�GJ���������J��H^p�� �i*�5�y���V������E�K�/�D&؀���-WP���,j� Hem���-`B@)~�J�m�cKD���A ���hQ�,?��<�����N*?-J.���6�@0��9%Q ~�;V�01�9�AM����M�E�<xE ���#���6�ƃ��ٝ�c��|(���l�
$�;rR�+�FB*�7(FΡ�`c����/A�:R,x�索�[�<�U#�E�9�Oѫ%�d�޹��`#e�˄.*��Nh�*vJU �(�8�	Ss�F�%�B��9���&�U"�)i�;�)r���9,)�Li3 Q�1�D?n�����.�d̴-hn���$2�S�&M�u4f�RPb'�9��� �b�.K�XNM�Q�M��D� 9_=L�?&{T���(�$��G�������&ڑI>U��������7)@!����B��J�����I�;��`-U�����7d��z��+�:>;4H@2%f@�uT�3���P\��Mn=��d�C(9ɵ��^ϒQ7)sPn)�I�i����}�ɪ(�	"/��@��~�C+]/����0+Г����2���=J0���Y�KY�MH	�`�b��`˄Zb*A� V?�>�����A��WKf5v�P���AjC�O���F
��YܶU��r�QA)�%|�$Cio����oZi�*��JH��g��ǀ(-�3P�����2P�����x�|����7i{�_1��O���7�/�wPl�^:��u7�;�0�_��}��M�A�G��#�1�N�>��3�Ǉ�� E�fЯ��tm�ew���߻1�M���ϫ�=~���Z���\ؐݕ���7�	ۋF����,B�����H��R����-��Ϻ�"��4gZ�p�C�*;���n�J�������|r,�MW=r���t�:�����^s/}����b���^Y�໤�?>Vx=���H���w��qhd,z��99�#�0��4���&bF9�)}h";Ť����&���MM���zw+u�9�gd6#���>���`��W�v/n0V�ue��Bk�SA����M͹x$!P��b~��^:��k1������|��U���3̀s/�=�lptk�� �<LRA͆��z�@O�Fx�[�0Y�+�uf`Nfq�h�!�����ạ��L�����v��<2�yC�MdyM��埄� 3k��({�e9��y���A�L���p�ށ���h"�ہA��qz�������uy[�"��p���}N�����?!dס���i�6��"K��5	�����Ύyuq�#��|߻v���d�=f��^�E=��i��=wZ�>8�BD�3��
�h����ܖ{|�����]�yN�Ʋ�dc��0�/$���3CYΝ}�A`���W���c�o&(Y�3�`�CH�5�u��nq�;��uWgS_��N�v�AO�o3�.��];��1�N����s�yMvU�!	�δ�Wi��(�ݽA}�K��w����]G�W�ۜ��j�v�%�y�v��g�٨��B�^,��}� �*�C�����J�<�s�MmD/����X�a�]������%Lw�%��?�k���"����K�^q���I����NB�kVS9�<��*f���OgԼ���;{v	"Ƕ�.�)��^X�'�;�#MR�:2߮��FQ#�W8tT�����i�c*,>xԄ�}2g���A2^42`1o}VnL3-�Pz�T�ޘjSz�M�!ֵ�B�gz|�te�;�X�wZyg�u�G��/L;;žN�q�ʄ�^�yk`'|���\kH�`���(�@�r�K)ʚ�o3�����gSI,y���8<��1�.��̵�.�ņ��X6V��?B(�&�|�I�Ze���+i4ٷb��w%fa�	y�����LX���Z��obZ����GK�:�ub"�EKtby��y�$ƙX��fc�Q���5��^��#q|�������-烹����-�_���#@��{�<G"]��t��_g�n% ��#U���!�uq�;�oU����ef��Ǵ��b,�&���SE����{��ȡ@��l��a�{�2�"�Q)��.=0;[�Xa�1��A1����ഋ�/��������vl�f@�#ȗqeo�?>S�G5� 8O�&�+i����m��um�R;�<y���Ef#����1����&�����F�q�9��]MC~ا���<�1�Aj�Y?��EDlB�SNѰu�(����3ZɎ֟4֪h�&�c�ը�ڪ}e����ȃ�	�����_)��l\5�CǸ�F?�u^X���z�xқ���q�՛'������.�S�j��7W���o��?�ʚn����nO�k�*��؞
��>���2��h���C?��vw׵��N\�f;���Y�3ߨ�	ƾǪ� n��6u섕�M7���,�"�3U%�Jd����j����a�Õ��egKO�ߊ��S�ʟ_��V�*�R��C��j<��U�Q� 7`�����^x�+�g#���bS����r���îE@;�{v�	������t�~��.)^���1ݝxS)0Z�]� �&�����;2����u��H1}�)�tSSV�˛�/B]�hC�*eL�zFn~O����F���-;�Z~����`I@�˃��w`ףiF�(��ԥR؅U)�7��j�����}�9�V��Av�"HDxt�5���PK   Th�Y��:$  �  /   images/f2ef8506-1b6f-4eaa-8cf6-e59ae15d09b8.png�Rw4\����F�d�.z��G	1zѢΌN�D-Z��NDb��� Q�%!����~�]���-޳�9�}�����g�'��XL�B  ����  ���'^#�0: �ejh��	��`�}t�_]]������9x�Y8\]]�r�f���4�4b��$ R��vNU5M?***.zz��h���p� ��]��@�BI]ORR��>����������c�蒈��Nϡ�f��G"ɦ#�S����L���cT|#>aǃ���v5"��~�W?m�~�O�E��/��u3ۅ]^��>;<?ܰ��bw�\��p0W�J��H�o$�t�7�=ў������(�ކ���o��􈸆s;��F>OG� �c�9�a��rH/��Kj�ğ_���}��wpq�{q��h���iŗ�D�Obsm\l&�9&���Dty���|��|���Ά��1�n�.��N�fV7�J�F�w7��V���D?A� �⣡����ۏ߼?��X�NmKh��K�Aq��9[i��-�����n���9�ds��R�Ub��W��D$u�@��`e��!��,��$F?0��)�����y�}�Ϫ�B2��<�E�T�~jH�C�yrv�22�8<�^�I)�=��Z�~��4V����"f�5��"�44��q�^d�J��K�FP����0$R�������ܛ����Fwm�Qh�f�������1[�#z�����T�4A���Ѵ{ce--%�N^��]��
��	qE�um@- �8b��a�����6���*�GG�n����5z�KX�`6�5�򚦦�z��X�	ɂϗ>���ߖ�����C���c�,�[��ˠ�'���
�vB�p�N�({����!�ϻ:���3��
.�|�*�^�!�	�UĘ�TrY>�0F����<~�:H3˂+���9T��7�
������m�:	��&�� ��O����$00�L�����f\���`���Z+��tJ__E �-'\��9X�i���ou���d���G�9����c���ji��8k�-j�]�i��'�].)��N�Dd��ݛz�y�Zj7�+�k�Rk��3d%�]@+�O~�mM"h�9Nˠ�uy\��x�<m�q�`xb�gfM���"�"�����o�PF�
矎�BsL���q�|F���D��J�n��Q�`�'s�u]�̞4d�FȤD;�ݼXx�c;��^�_Ur���6��T��>��0Z.˝T�ׄ�}�K~RU!��L�p#�q�uU'�_����G�S�?�����,�&⩣��t�L�N���lܩ9D։F����Ґ�wg?̢o�� KF�N�s'#-��t�,ڣ���W�3�뼼/�С\�Oڨ�,��(���ɑ�׫��9u�0#=��a&D<��w�;etp�ྠe�ǌȏ=��� �Pi9;�1*���Z���s0j:�����L3���Yvn	R��Q�Y��|R�cڄ�fsA��_z���?ș���g{�Ap/fҒ��aV�R
��l+���杲��g�u/�3;����{YG�Iaw�@^�}�hLi� }H��}v���^�J�GN2!���Jx�sD�r�~����N1����H��J���ߓ������R�7;�R��+��!P�<g��7�C<z�=ILgY&o�(��1���uV��^O�:}�s�Bv��2aТ�a�k�&�����|�iA6���Y������*�sY��h=+b�A>.pRD���U@�X[�X	�X���v�E<�w.W'Έ���n�0����Q�y��N߳����Eujտ;�y:��D�X��y;�������?�MQYe�]#�����Wp@!�o�ʹ�5X�6��gF�?�~�ef:��s�Sj�p�'k��Bhdn�J��O�����-�U
����� �\�D5�9y���g�W�[����l��8P�2�)B��)�~nr��)������j��c�̺/u�����+�Yꪔ�2�d�0�r��K���F�����!7'��
l��Ű�ke�������M4䝥��/���5�a��k�7�nS��\��ot���|e�#��F�
^��teB����˰�U�|��� ���4�:���Y������٥�&r�hJ�k<Ǆ�*��d�jl��?��^�Fs�����(	�r�jvZJ,<gc�фl�I��R_V�{�|j��nT�Idtyoia����@
G�+�{�SW%�W�'��9��������UFe��9��s��ن��/7�Ԗ�����ݲ���\6|�����j�g]��6T���ʷ�C*��:2�f��@���Y�D;j�T�L�+�ϺAn#�T\��r3또7�3���F�3T��އ���*��̺���;�R���/2@�[�-2�o����[Xr�	A�������Ϝ��S�tN��)+�6�a����?B�V�Ԫ�p\ƄO�K��\6W�o��ݘi�����uP���a���a�[�F��c}&O���r��#���̠�w�5g�����z�R�}�#�]�
��=11-+��׫�v:�213��7�k�������JX�  G����ch�é��i���O�U�'y�{��m��RX�(�κEs����u��������Ϧv�+�ۂ��9݊]�\!1x\��x6w�|b𜸒��o>>[zA����)��$}Kp�Cˤ�MӬ !�y�a(��~i ���+DQ��B-�Pi�1�f^s@@�R߉ai�7�/��9�8z[�S��ž�N,� ͠<2�uj�����%�h)�n���@�'_�dh�KD�һh$ɍo�A���7yF��`�҃%�O�u}u�.D�+���/$E+M���vy�u�П�5u�l��7U�s���_�P��o�V�>�l���,�O$�e �@���\�ދX>�ejS���k	1ob'B��ɕ�K��lqʐ'�&E��#��|�X��}C��9�̺�`�Y�n��� �NK����y�Y�ǖb��4��D��B���\4w^O�;��Wͮ��q5.�^FqF�^�=�'e% �G& ͹�zt��9���&�("J��@���(��Z@���%�����(��{g�4�ء]��ν(��M����e 9��������;�[�ù�U*3�������݅V��Qo`���&8���S��Q��^���n��y��m��a�.��&��bl���A$U�Il�
B��x�݈�2g9p�I��;��F?�����������=6R��V��|i����fj��@ܛU�C�,�,x�3�	$&Kq�6�������jL����5>�&�ŀR­��_a	��?�o��r=H~z�qY�����d������EH���)D��g�]�tb�;�W-�ut�ni:^&�R],��4ܸ������
�������	,8(�d�~)R���dcg���] P��9H��|:����
��c0��Bx�
�&v1��_ʪ#=����G��I��U��?�J���"9����"b�ҝC�C�?ة��O��n��%�52e�S��s��W�*�e��˴,�����{A��R̙��������s����:�zi�R�!��e�T�Z,#p�s6/E
WW׽���Q���T��7����JFdF�=ߓk 2n�bV$䩎<|�oQ��� ���a�~����'�|��Ҹ��2)n�jA��s�Bl9wZ-i�|� |�QPNJ��X��p1��ד/�4�"C|1z���
"nN�%��*�a��H0_��D2W���4���Ѡ�Cκ�@V��0��y�`�8u�o|w�UFG��J̀o�k��n	=�o�b��PlW�xG Hw[ߠE<�`��O����cQ�n��F#��$hY:46/q>��qv���K��.����
�������Ux�K�(��*��!h��=K���Ld���o��8�Abٸ�e%$\(��5cu�	�H3���$Ș��z�{yH�%�u	�:�01�NG �9��1�������������-W���0��1��wc���i�ꇅ���������d����`��_Y�@b��K�G�J"�|�L��� ��Sr�������p�\M����W��$	�)eN�GVF������/���Ͽ4�:B3��!�����0��O��#�n�������to�*'I�g�/t��� ���{S%�6k�&\4/#E��X.��C0�S���n`p@�c���b!�hws=�*��dW�[�{�~H�H���e�q�i���aw�
f-w�7p$�a1��t�@����ӆ
�Ә8Y�ew
W��n:ʫ�ȥ�!�eu%JK�z�5�����w�G����f�EA�T���㻕��^�����	,�ڏ�t%}qdfN�1�u�38(�'"�ZV����=�P��I *H|0��Q)����s�Nk�S.��P�˸+�q��67�i������GM��p�Mb�	��/�-+W������n-c"�
�-�J��G�[��CzB�1��\(�"�j�Yh��2N�赺,%���j''~�"ʵodz�<It^��@ް��	���z�U�=52R�W��w�A��IgQ�w�:���*k	P����p�w�T�?<`���~a����̈!�B':��%	�,����+i����(�9K��w��7F,��N�'ެ���+��D0���_�Gs�>�>�?���msF.џK5^[��żV��r��v҈f��\��R�yf_������T��2\e��&�l�wPf�^ֆ���Ly?�4���f�Z_
]�����GD��^������`��Tn�
lL�,���t�.�n�3�*��2�
�1��˄�:���"��ͩ�>� �x1}7)�}$�d�%BL�ףQM7�{Mgk�q���:T���'���Fś���c���I1^x̟ov�(�]�|�z��X���F�*�F߉���Ί��$�9�W�U�GY��o!I������\3���ŷ���֛6ݜD��<1��x�W��	%j1"S�r���ZYߒ�=��Q�~�0��8�b%�&�*�L�������f_g��w�N�a�o�=
K���?�&a5=b�2.�^�(��V>�X��u,z�����:_�uuZm���0l%�x�c!�ݹ0����)���o盜MJ
S�N=,H��0PZ�І.������T���J�Wt.��}\Cg	�+�'�X+��b /�D�l3�Y�b�[��nG�ʐO\�Ph�V�/���b:gP]�w�ߡ�KC :¦
G��P���:���nzAMQ�mw�{;��" �͓T�nܒ6i:���J�v��A�eO�F&��v���tS��ֳ�S��ט`R�*�n#��\����+�PD�.�f�fr�9�9]��F�*t�/�zջ�����HG1T}%i��K�b���	K�P|��r�}��0��;�-��@D �X4���W��l��	e��4lr�$�A��$%�Jv#�,��՞�}lJc�+�!Xt(�UeEjӚ�[���^�Y�#��� ��`S�J��b�L'}.O%��H(��9&��y+�i����!�jy���F,WlR�Gg$�������tҲ?�nʔn��yFX.aF���f�:jW���0�NPX�k��s���'��`C����o�ҥ�^��@!zY5~%s�"`.���,�Ӑ/q�R͢�����ݰ�N9)�ˢ��O�<��g��
��A�b�z1�N�+�[p{���)1�Q���zxI@���c���pzJBvw��6�ʮ=���{q2�/~mH\Zo=aAÎ$T��Q�z��$��P��r�>��1Ta}�K�������jF�Rs^U�L���DE�]��؋"n.��}pr��}�ܨPm6���6���`N+`+4�)������W�R�MI�d(RW_胓��N5N�)}v+�A�h�hm.�/E�Q�Nr�=�=o��\(I��@�G�ͫ��L�$a��:��G<�43�.j�ɪ"�ũ�%M��M�B�g����F1ܝ���&5Y��sA�#���س<��ݔ���L�	lba���P)�\O�{X�c}�g	eqТL��Q�f�.
�f�l$p}�k�j�Q�PK   �f�Y8�w���  ��  /   images/fd1e7351-dbfe-4fec-861d-4a74217661c3.pngt�eT]ݒ6�qww���=����7���N$xpw���!���s�����������%O�ڟ�eP	A ����*�A���#���'@��,��)F��A\R&�	ܥ��՜,ݽL\-@^^^,6�vnf&�,N�V'�� 9HNRL�;�軗7��@G��#WX���&$2RU=
�(�h�OLR���
	B�X�*�>�z�hP��2���H���;�G/��Ga�������0UD#�� �|y)_k%�E�	n!|�Q�xH��:o�'
�󊳡k���AV��Ehl�atܽ�V�}�-£�z��4*�����R��[C��sN,�4����t�P��P1�s��k�a��[��9Uӳ��$ceoZ���Hd��nD�N���z]`bX��;��n>��v���*/2��Ю+D�Ѕf2g��
ZU#��*�*�Ɏ�$�r\�gq+�R]�P��blz��r"�V�m�BO���N�J�Ӕ1>��Ptǟ��.�;���r84(#!*&S�����C�,�g�"��oá�l�mI�b��k�}�*[�:���rF�չ&�!O1ogX���@*�n��^i���KtW�U�,�p��d��v+�)tpʊ��мb�!�2�L��uh<�V?y�M P��<�	���?Sby�J������Hb��<խ:9�c��Qv|З�͉�c
�:���9�	�(���)HBOT�����p-��b��A�Aa���b��HȣqH�_�ۃ�#J��s�'��L�	B�r6���ul4{��x��i����=8�O�\QF	A�|�&�
>�9�Kv�mb�U��tbDev;ORq�`�o�Y����v�G�P��ˡ���h�3irq2��[�&�����l ��E�lP�骟Mߑ�J��2��E���b�RE��/��m�*�t�jz�Ƞ�*�M�'.a�+F0�6@��.g,S�P�xZ ^rߍ�!*���,�)e�q}	�z�"y�L�bTtE�Bs��$g.������u⾂)c���.ȉ@�F���t�>�b�XC��433�024rQ�I��ʑ��������H���L8�X�o\�8�qgt�w�t��|h7��*�� 	�O���bcP�����?y$S�>���Gb�gT2R��dܕ�u��|F�S`��Gz��)K�jY^��2��Fl������\���o\��8�\G�!�1&h�A�����m�"5��#��
�A��x���+n�<X~&Aڷ�cQ���V!'�졅��rx��}�Elv�4{↽) ����o+~i��K�#\�o�XF#��`�kL����0�TO-�;����"�Ck�������G�f����`b/ ��M��vgC�1|���Ou+�����ܕ�+nR�Q�1�.��7 f ��̫Č_��zE�E7�bc��v�ɑ�*�j	n�g�_&8s�S�J\Y`4`��J����g5%e����5�
D�6'9�eS!�G0���s��s�~�ԗd*@���%	� �[��J���0��)�nV���ݪ4UY$���G��6)���Tư�:�&�X?Ƌ�j����^�bs�7ߺ
J�M�i�S�ZV�:h�+zO�8�֕e�8DlF0�}G�SM.=4)r�1Mw�7��S2��Hb��)UG��>b#
��+0�B��6ϸ�������Y���Q�I��F�b�O��&�Y#
忶�&�A4Պ�@퉲��%�̇���5(b���(����7_�,�r��w[|�6�.$��W["3-��������'27DMbɥGg"yS�&�A(�3`qe�Qѩ�,?��ol
�Mb�KN�P�B��L�V���]Y �@�q"׬���p� �Lg�6gn�::$���/n�(��SʒĴ42��FE}VXD) QJ�|� �7�J&tQ��F>m�wzȥgg"��$�C�5	�:4iF��6/�$r��H{��3p�H�M���T���n^���ռ3 ��'C�h��GT�`�i��m�C
F7�;�V�~_f���BV�?�䪜B9����[�Ҝ������B�t���a܅�oV�ҷqi�t���a؅�%۬��/Z�-����:�B��/�֨�`q�{`9���@��"�k꿚��]�w�����C��0����$F��}�I����·�T��Qs�6M�C1��sX�n��V ��M��Bz�5���&�"\�/}Oto��#�ŋo�x4�3SHI��oWC=�/��@p�r�5�4�{f:�Yᖧ�d"�r4+���({I� | �B �!�{8��;�>��X�@;��Z,��l�qp�.����+����VR&���T�vL�Ц�ۅ���N�<��ٗOt^|g@������s�<�
�K�\�*���VT&�̿��,�F�ㆹ�-�P��4���:��Hy��e�=��f��Y���Vκ�f[j�!�Y<�&�}�R��u�r������V�v�Rݩ�����Ue�Yeu �d�R�{g`���y.�ddd��H��=�s����=q8���^�"l,��R���FJ�@?m��a\��-a*��T*ӛոe�:���:�
p�Z��A�f��T�]Hj�b���T@��1 �ah�i�d"�������3��h����_�|x���o��D�_�Ə��*>KR��뱖CJ�$2��v��fX�4�S}�Q:Q��:pEsR�#c\M�5�2k�̰�CK���������m|+'�dQ���^�(�r";E����;:���E�8j{�4Qsz $M�G�j�@�ä9�ˬ�Y	�׵�w��z�׾���>��h���;�Y'�(ݕ�Q�1gJ���,7f�O��g<C.��$d�� OǋG������Rl���f\m)ts�F��O���s��֥8=�҆�w6 ���]s�6���>�<|h�^��>�R�7.`(��a���gf\�����Rl"�V�D�J��Qh�1�<��֊̰Je��8��1�f��<�mUEH�'W�]er�X�A��hv���N��B9��vWC��i���N�12�X*�f�J���.�����ԩ+��N�cN+��KG#î�t���%��5T�����?�t�$CW�n	(��-�z�L�OѼ.��ƕ1�������(�Q^(}��v��I���(/�-c- 9�?y�]��ha?�R���+3����'�>ﰸ���d���z�a����^=�,�k� AP �W,��:O�7dcrP��8.^j�9>2lh�1�/	x����V
ퟛM�J�����.}񈌓�A"� �0Ɂ�^��U�3z���s������
�7���L������.CF���*�Ġ�Vc�儬vݔsZ��R$�2����`��3� g�)��� 敜�[�����^�3�<AL�J��r�ވG�G�>Ձ�ߴ���l)O�mJҷ,��v� >�z.Fe[$o�s<�F�,�xL��̾����}}��6�q	5����%��1��ŵ�4���=�HB��^%�m�������ԫ��~��ch5�՛�%��YCY펈��X���]�łM�&�"$�,��?�E��.����)��V���4R�\�nӱ�N���l��Nz�h77DȚ�����>9ѫ��߹���F��|�Q���ex!��z*�=
$��_� �y�tʹ�ǈ�Q�L	y�T�sNi�9��Ґ� �yM�7��)O;���)�̲�߽(&'�������W��;f�����=�`A�ivj�=KAͻ5����t���-P�G�:d�f`,��y��Wߞ�U l�x�;Eؗ��`c��(�q�ÕL������Cp5�7��q�E���4�e��F�R��P7�ݚ!U�h�Zz�c�����\���c��?v�cm|��������b^�_�zG��_���5泩�][5��q�J�.VVˣ��A��Q�~F���5��������+�,y/�N;�C1�XSLf/&�&�}��E���V��`��ow6wn��vj��ߚ̳ 8���[O���lԼ_F�%m�[y�U\��K/�u��FXAξ�S�^��xA��F��;��Ki�M�[U��۸#��j�$�mE=ul���Ҏjg�2hɶ�cA�%��eO���ǒg ��Ӂg�����U��մ�*�^U,�3g�{i��b�[����CvR3)��,��r{��i�S��'2�'�Q���R�>��j߻]��
���9((�=7�g�'�¾�V���BJ`^���#�J	-$Xy���	8S�wM��d�0��z�K��}�d+S��}xd�&��mH���@�0.�6�-ǭ��5�1G-,g@��s�boF��g��.����*D��+�A��P:�a�״f.��f���i0�!����J4�BM����JZ��)��?Ի� >f1ev���؜	R��؅l'=JD�6�lFnT��`�oщv#Y"#em�>���ə�*�
��UM_�_�2�pSC�Sx0��*68�]54_��� ��T�V����V���:�>���&L_�Ru��0�,�Ϩb����k�Բ�u�w-���X���Q���l�?T��S�bQ1#.�u�m���@�T����|�9��7v�ޣ2�P	���_X�/�R�j"�O��Q�����A�k�	)i�gR���]
�%?L�{��g���v�x����ZT�!5�%+��ɿ8�Z�~��"E�UW��$ ��+ʊ1�tw�X '�A�=�b�B�Uٌ���xl.a������|0	���	��G/S"kCax@��8�*�c���C|��	�z��7�7����� .�M����׽/w.�}�$���U�y)��>��US�PV�js��qe�dy��yo��<���L��F��E��|Yj<Z�b�z���0o*��O�Ƀ�4P;�v)�֒r��FTIw��y#�s2�6�N���"c��]ψy#ɟ���b���٢/"�l���۸����IS�0����a:?��B&)bl�M�<��pT?G=)Z���#����Ŷ��4ۍ�l;tXW~L�/7��볝�ϩ��t��_�"c; �������«�_~�_#�k��&+���>Be+�o�!mX�rX���x��hޔu)���2�B��H�ĭ�g�uë����j`��R�X+m��צ[�ւVǫ��:<�p���gtU_�(䋎��pP����}nMIj��?��L�A��n�?85�2�?�#��WQ1:��C&1�28j$�{tx�%&��\�8fvW�<�)$�S����:������?��S�h��#mx%�s���W��9�K�w�j���m�*�� J2R��vx!��!]���#敗�緵�Ƿ�����}W��o�!�#�x��/$�eX�-{H"�UܯAJh���<��hEq��;��OA~�]��0��ĢB'$9��j1��h}d��8���3���šg�:�c��W��[�A�$����}��]�����d��_?��"�o��O�y[�C�0�������Q���+�^ppMu`��7� hH��������������+����J�ץ!����M��'��H��S��?Kϐǻ���gI�1�kՋ���B�b�u�8�4R݈q����#HM75��Z���M7w��F�5���͌Q��^r��׫	�m�v�i���93�Ot���_��.��ٟ��.����8W��[�ǘ��(W�Df
��R�Ո�gL"C��v+�Iv���Ý�x"�{H;��l��9����R���`��ߩ�N��y|o^��ؓ�EҪ:�+�#��ɶ�
��*�K��Q;��8�1x��YU��B^¹���yR�a�BA��/o9��MqxW���>�@}:T	E��M��n�&��V:���g�_l�|0Q��m*�n�&���2���mSeR�&�cx�z����	���6�Tx�S��i��=���?������O
�bc��0�\8���L�"�ˋ�n3���t�O�,H�e�H@~W}͏��P��V�+�T`xr)�TOLb����T\���1 HWQ��ʃ}��ԫ�ŝx�1����y?|'x��.���٨�+�P���z1.�����>*L�,쯅�$~��"]O��N$���p��u����"NF5{�Q�m�O������MI����j�d>�u$9��|g� �h	�}����,-�\m���\ѦqV���M����/���7n'J)��Ts�w!�S�5��aE���\Yr��*�<�'O11�Pc&��ߜ�
K����Ǝ~��NB������Q�����@uf[߿�W.�`���Z�⤀�L$:����m��O���|o��{Ԣ�""8ȃi�M���á���wm������c����䚩��;�tr�e�Į��T�q���6I'� �4�u����2 W�rY rSin�����_9E0���4J���	v�'\5��N�ˠ�*�3(�� �Tߵq7F����B�'^-��3��������ej��RSv� ��>���o�M#1���|#.xmon��0=�3F��:�PE&��^BM~�������T7�&�fWr/9/�1�m������e�`YK� �.�k���0��]�+�#0a��V2�ZBh����#�cO��U���#!N�`¨�Tu������]Sܽ��K]Y��#�7�?N$��?����W�IT&Ҡ��63�j�yn)���$}�><熶u�ߚ���T��.���;7!U�
c90\��mx�.IM-�g��k1��w�v��7e�[��TL:�����!�+:��i3���8`�f��M&�VH 3�[�d��$}̯�"�, ��#w�ϔ�?�bcqo�)�QL�6�2��3���jԂ?�vk�i֦��ja�IM��qb������(�$P�N���Ŧ�J�w��M5�-p����?�Wd�C�o*����ȝ%��3�TjJ��f|5�m��,�T�w+X|x� W7���*�C����N.�8
T4��}�T��	����6�+yg����f�z��T�/���*F-zj��&sU��/��3I,/��)v!�|�ĺ�t�=�47�bj����k��4wv�H[9<�1�ރm/<�R`���T`S��c����b�3�����L��4�	5-��D��� �e�w+z=��	�N%!���N����j��%�r��O>N���8?�)��I,?3�d����K��j��J#�<4�b�h���L~��S
��\��v��
-/<=`4��i��7<l�*ڨ"R�,�r�UFU���n#Ü���k��;�D<��A�����j��} e\@��Ж�R�����Sh�lzU ��t�jv�ۓS&'�V���d.�	0��ߋ�o���}�H�c��ešA���i�U�����C?O'�ԑ�Lp������r+�P��5b3��g��zz���5~b���`���q���I9q�}
l��J0�L�r]E�1�c��᪓��?�=��o�OzU��s£�NG�v1\D"6E:���a�^X����D5hU��W��L��s�DV`�0�r��-p�g1�H{�@��]t���T�� 2U����5(gd@����K�*iL\}G�"����pQ�2l��+}&�Z���9lݠ���ʑD�|�Uҁ��[bed��Q��Y{ű<O �FU�:��	�?���c?��T��*�h�,I�@$7�'�eɪ�$�XL5H�����2	h�8��?n����o���Lf(�o��0�i�8�pK�^�����ȑ��sa$�B�;�?s�*A⃗�,����ݓV@څ[�(�!��wJ��|ğ����3���o�6Y�e��&���cp}��~�#����?ҵ�"�&�*��fETО}��tխ�Dq�Se!=��M2[ĉ�����k��]��y��64�Y뱱�p����������3��A��f&�\�$J�YOW_]��#��ʏ�t�)�s��3}�-��eHM�]�?�-��fkOn�M�J09���J�i9*���Y%�"��䵂ڙ�w��@wf�A|��x����j�H�rn�j[*�q�l���#jzS�B_��U���T,w��`�OM�ٻN��pC�C���	I:�*�,b���:Y� �C��<��PQV�=a��|'�<�B��.e�����a%�i��2w��]o���>�{�S��u�3�1�Nc���){��把g7�p���̑�	�B������Kc�����2�ʵ��v��[��'vz�#Ó���}8DÚ�k�z�1�ᰐ����Yko#nc��L���I���%�����h�v�B,5X���%���T:Ɗ���H�u�����p������!��r%H��c}�x`s�h|���ߓ��\*ɰ���Jl+��c�@
�|�z��f���-�&��]�i[L�!���`	���q�yrb��㘰�Q�C::����r���l*�!%geЧ5�f��O�=�;�mC�ެ����S_M�J2�����(�k�#�Ō���t�3�%��e�WG��
<�W��_U�s������c�k�.�)��'m���n`0��U���i`���/Nmp{?��g��no�t��\� Ǩ�F0����x�B8�O�B7;!&Nx3���1��
��>�U7�R�K�����R5��w��~>�%_��`�G���(z�m/-��pC@%��ij�H����$�E��OFH4Xj�J���A$���k~$�e�}&|3.�G��ʺ5?d_�{��z� �<����z$�\-�si)s�`v6_C�p���]^-8��h��yzv��{�[e��aq}���:�wvgW��m~�?l�do���ZN�]�ϝ/}�x�����ڵdM�m%�H:�7ܵq)h�MVk�>�{��t꽼�\"s.(%WLjU�j�֥VW�e@�K�9ޙ}��'�	f�|���-����͍���(�Z�s(�r�ӼA�D�����56v��9Ͻ�YMڈ�-@h��=�(K��$|!����]ܗ�ά����n&Ґ�`�I��~R��I3�ý�j�'^N��,��E���ƞ�I(����	"��� ??�����v8	-81�/�̎M�sj�,p�.���d���O��亜�D8f�����fM� O,�� �GAUϓ���4�2�0:���b�`�q��]O���]�Y��`� �E8�{��S��Yy5��l��e�)Q�I�։���3��+�b�{�����3��fx`lltY/�A���������zW�w~�Y=hn:��፛?�b~d<��:��S��u3U�m�U��G���������A��h�� +�~��*�F��4 ����J5'!������ta������yn�
e
�0��62�W?t�oQ.ѱV@Vn,?*+�c	�s��T)i	�����"P �{�-ݜ�c5e��F��{Z��mﻡ���
���ۀ L;L:O���}b���oa���{j�ߝ� ����dtB���eѼn7��pM�5�����{���Hd���l(��`�A��LBQMD�F|�iw���i��-�b]��͂��p��P�nY@���cT_�.Ywo�������jID�bh�y�Q((��}����h���}��� !Gۈ@�ȁV���C�p�0πɽմ��j��{�[�Ht�m4oJ lŘ�Ǽ�T�?�*^[de%y>ɐdS;&�'M�����t �W/ט~R�~�k��%�؛̓BDT�l{U�<�[��%�����i_ߩl
��B��E����zi8=kY�v��$�K���|ۙ#2���dɳ��i����@���;��� [L3À
��&��ۆt��5%�e����c�~ N<T�9y�Vo=+X��Ei���g#���\�d�9��Čp3�ݦp}e�3��>}Zy�N��z2f�m�c�~��aF�>KȌ��;�Κ�̘ؼ����c`H�ҙ8d��	������e����x�#�l�C`6�Ҟ���mWge���Z�CPu>ts���R�%��Ȧc��]�W��==��k��0X[=׮ߓ��N�|��+�^b ���o�Z_G)�3W��j�92�l{(詭��y:����n<���&{M��acpxHBE� �P*�&�����gO����q�%9D�Σ��
^:�1���,e?���LwCM][��iwD�v1<r53�$u>��BU�ҿ��_'�$\�R5�9�v5�7;}w;�m {���[���G{��nD��-���l�^6�:nj��ã��7�=��[�݈��ib�IERCٱJO�&�۩�.�4�-H&?��7RK�-����w�Ԓ�c�����(B��̯"��
�������Aۙ�0��먝���gdЊo�	�˪��U����z�·����c� �_\�k���c�-�2VpC��e
zo0�����1Ds����s^��Og:��f�h/�[��xU6���#���޼��ɞD�-'/H�\��a�l���}I� �G&�j�t�sK��g�bW��\#�=�� ei�΍��4���� Ʋ����VI(����u�f.	����I�����k}���ʅ��-�v�:��I�Ѯ����<����x�=�鰘#�����l���6�js���T�i�N"��W{��j�h��+�ox��̻ C���)ѓs�E�pzx�͝]��q��J��͙��{j�a���j��+��l"��΄.��+�[��9��s�*����P���]��z�s���fu�t��'�ZY�5��/4m>��$�.ӎ��`���{'�ǋY~V�R؛�(��O&}��g����N���ڐ/6�v=f��(9Tl�rXQ��� }B>�9�6b�sd@%��� B���y2W=�.^�^Þb&�^ԫ���Y��ؗ"�h�ܪf7�I����d��l֕��t���?�3��8S�����Y�󭆊��x�^pNJ����1��Yǂ���1�:s~�������@�����h�a�b��%�zh�a2��hOzfl���G�e��ӟ�e&�58��Z� R%v����-���$�O�_T��s�M�e�>�{���{��Q�7��h�9 �>..*✕=�[j&d�7bz\x��P��r$�Y������Ck�7ڌ��>uK��d��|�6�ǯ���������q��L����9Z����q�j[��6�.BZ6�_��\�� 0�콳6�������;�|�J������}y̞ޜ���ޟ����t
����Vj��'a�׈�BW����=�@|k9�4�W�G�,q��n��~ӺM@���~}v�EY�΁@�U����B��ŭ�AY��―��=�Ps}��V�m�E�3�����H@�����S~~˄�4��|u�խ��-�����Q7�L�fTE\�|9������� �*˻N�@�)��
�|�+˔��x���P�M���\��������6Na;���ĵ@$b���d��q�7n}��1�^���cBW�y�=�_�^絶����*���q������� ��ǣ�]x�� �҉��Z�>kN����2V��%z��d�t�󅹌���Y�ـd��<؍//�Z���A���v;�>-fUy���yz+��ܾo��sK3*���/�&Z<6�S4:�s�U�V;�����<�J(&MF�'_��n�&׋�ʭ@��?i6�������nk 2�֤�b3�>��
\P�\�=~������>�DG;X���O{E>_ �
�UV��@j�m�A�����p7-�������GY�q��^
���?�n/�\Q��Y���ڒ���|i�"C����/� k�C�6" 
���9�N򕡕	�8��IZ�x�iO��G��0gD���
@ț��޷@����^h����B�o���v����S&����!h�]�" �4i ,[ϐ�����{Y�qc�&[BA�2X��8�x{�!<H�'�zά�G
 4�;�r����� 5ҷϘ�4��j<y$�ueB�w��P�ԍ�p!&���ߓ�<Jb��^��R�ޏ'l��P��h�-'-�)�8]M �L4���ͬ
��?u�b+��q���o�̑-nAy�K#5S�a,�ˁD���鱃7Y��[�=��Lޯ��ָ��h���L����ۑ&q�}�[݄ɞ�Qvv<T��n^��&JF|�r����H�����Wr�;�h|��"}EH"r&�0H4�L~\����
��.�E,��v�_<��9�B�Q�8����J_~%�P�n�h��l��e�����gN�,ը�
�����.��w�����5&s~��P�P1{�7^�D�v�����P)����C$�������:R�6z5$<��!�~$�����h���[S��y���Upm�JI\��k�6�f��A�Ɵ���vF<�?��;�q7L�]�M�1��b�R������ŝk��V3���WR/旘��Ɍ`�jQ��J:�t�$A��[�8�=��<����Dc�z4:���O�P���t�/�>�.�ߜJ�ޕ�:��1�d
�i�a�,�����3�7�8jH{�,��.��=�v�GY�-{�ޏ���~n��5��ΠMN �4��z1=o���m�ZG�.�l�An�[������`�!v��� t�0P޶y������{|;n�
v�E~#�����-���4��[�?IO\�X��t��S�����\p��oHa�t5�b-Էd�u��U�:"�4�>�t0'�Glǭp����<���r-�چ�p4}�<a!��a�|yFu|��K��N��z�  ��n����>:Z�ĥ���b�M9����BL�\�������#�~ �i]���]8�ݏ�:r{��y�eN`f3{#ާ+���k!����U&�Lа}Z·:�5?Q0HqÞ#ޗ�o!�]FU��8�5��w�TqKq_}�	c	I�|R�D��&��_�l৕/���Om��w;d��0�wfKb�����y�(�(u��\��u���Fa�������L�A�\�_��jP�bPihX����k�!��I�y�eA�9�f[j�3%�_����M�T?u�>��ru���c}/:Bz��Q��υ3��=�4�d�g��0&��?�>m���FȌ2[b���6��6`���(����^8��#���l������۬��&__d�s��_��ӎ�٘*���oI��8M��,����i$�5#�#�� �c��,��|A����2Oӟ�&�'�6��,s���z�����/;�G���.�Y-d�}VHYݍ�Pg�Id+q�Q
�}���3��J2��F:弜�z;�yVU��������.g>�u���@�;r���L����,�ɣ�DԏM�Z;��F��J�IXb���cS��ɍ7�*�RX������+�X��Y�_��a����������|xg��q�7�u�c�~C�eY����C
�]@҄7��p�5�4���]}��lɑ��
yv�\GG?��fz~��*�Ts��x�
���u�]�k�W��Fч�	�Q�������W��׷h+��M�hftK�3<���S����7��|!��~�y����bIc� �v�w��cb�����S�J������Q�������X�Сň��XI��퇇$�߼H���~� P(u��q�������T�L����9�dm�ë|fUr:Q�QX+d�^d$���B����QX)�q�G�+rrr�J��x��u/�}[��!iD���[���KQmt"�Xͣ|��5��]���~�^nc�u��l��c0J�o<�C�����E�k~	�o0嚱{E�>�L�Dp*:j0��_LE>�Fq�o�S��fKگV��ގ��yk����銀޷d,' ���!�
m�37�^�4�1��8;��]rfd�:̌X2�bo	u�H����E�C ����&�2�2�W�uE�J]��\i)I�av�|=#�Z���ݬF���1��Vxh8��{�l������ޘ���������p�����f��_�l�� ���znl���A��C�2&�V���7+��!����f���9\��M{����-����>D�"��[=Ku�@5�i�H���7�8L����:�۶0���/.��3:���fޓ�T�D��b�e��[���~\��S����%@�����͔!"����G%����$z�)bw&�v��'ۆ��7�i	�M�T���"����c��jD������LF�F��
�!�4�[t���͐�wFd�o�T6��s���~���f�Q�I�s�����M�
L	i�G�Gٿ�T��'��ʴ��~r��ƟLw\�)����\uN�@���G���M�s���	�̥�M������[M	]\Y��U��d�2�a��$qv�� �<ǁݑ��
hV�o��(H#^X�@T�d��kl��ZW\G���\�D���Q�>6
Ѣe|ǈ�R|Ȃiߓ�_�Y]>�h/��I.��ՙ>�p�g%�-�5 ����g_���&Uӿ�4�(�zs�A؄���ɉ�Vpj�E1���x3�p%1����鈯��vBʅ��F&U(\w��|6a��IhDI|��[�1Z��D��i��q��}]��ߝ,�T�y���ݾy�*�7�*��n�F@�������<���ε�*�22��$~��T��h�s�&]E�Vo(������{}��
��o_H��.O�] k����DhF?�n�YRq8�(vn����0?����`��ƅ�"o�̥��cx���E�Z]���l����@.dd�)M�c���D�L�k/�\�>"Qa��K?6|��q����ff�i�y��XC���Ijq���>�Sg~��hr����ř�N�f٫	ܛ�ݲ��~�1�#��p$�yؾȵ�s�����d5q�=�,���t���iyN��Nj��tL�/�ﶵ���ɉ�e'�����vn�,�·�_Y��s|���~���t���{n0�c�����ŢR:����݂w<L��*�i��\��t~'�>Y��f�aPꔴ^*Uk!��|4�����@�v��A?G
h �����ͣ51���/x�3�I��h�_����7�*V+t��]����F�v�:OLM�}e�$�����Fv.�͒�O�R�<���u�F��㖩��?���h�6.��"���vkR��5�JYhh�5E�W�6Z^���[��)�	�_~���3CB=��9�(5���������� ]<g���������v��8U˕�Ӵ��{�nӺ��o}���
�o5��a���� 2�]�E���5P��cl�n���S�6_!V�}�#��bi�j�h��Vԋ�Qo��8�0㓲��._n���7��aD����C��1���ɱfM7n��k��;].j�k���#2 4q��7ȃ�̝2gM���%�G}3o�C&³j���b����I�Jb�MkZ�i ~ g�>e(�����������ҙ�7/C�Yd�~Z(5�7Ii醆D�*�A����]��X%9�E�Q���w�[�q�WST�A%+�-��/t�b��I��������^�8��X���L�{���EX����`�>�1Y��$���? 8�M��gP�����{�#���"/h���NYn����7�W�$hu�z�KN�B��N��� Ѐ��,l���f�b����gkV��5ӟ4���O�pG��ø��s#�����>����.w|��Q�LBR7:���O�Mݽ)]o������k���s"�ΰ|1:��f2O^�����H4u�zGN_���p�����Z�^�?�x�b��������v��`�<�h]$�89��o����sf�
��2|�S�zE�����e$/p���`��g	�s�0R�ĳ�{q��Ӡ���,NA�����ޯ֓e.uǹ��*����{���_K���qG	�2���eT#��|��Q��N� �3��C�Ņ����[S���hi*��8��L�
e��R���T����sV��3����j�$m�`g�Veۺ��v�R?�<����C[�5x%���`ۊ�pq���"ph����in�/'�t����{0>�����AZ�V���L� d+�4eO��lԨ#��^"��܏�ZK�7�G4�����.5x�Ά5��b}ꁋE��`ShQgͨ���-j�&��v�`VC�+���J��z��9���"�� h��F��Ӷ��D)亢�3�q�$<݀�5D�x!"w
>��+�.�H;�h��/�����{oCۺ-U�縯�q]XX��Rk ����k�ފ�������D �`���.�x����m�%��x	��>�["���y�ǲ��LW*�I4���I��!��)f�� ��G�m@ze	��(ح)��tX��n�cNy��Ǎ4]�?��sH��E �#V��t�Jr��z�/b	b��c�B��;��w���$s=�~s��*U��Sc�����!i�5�����2�;���^.ߏP�Nz�yE��ゞ��=[�9$��y+�y>}7,�mw@^ͼg�����~{����������>xT�ݺ��#15��1�߃K$cv�"�q��O���zn�~�������v�/b}�3H{��]�N%�{5�}������4'ec�L�H+�8�����!u*���)��_�NM6[`!-c�FW_ 
>wH�n>��Xƴ�j��3A&<��CI�G����7 
��D�+:��~�p� �=���,���={��[����0�%N�|���Jj�O< �I�\'V<r��(�p�z���&~��S�e��N���*�xo�*�ǉ�wg5� {�ۏ�'�|�d�.�sc�q�Ƿl�����j���EAT�D���R�w��+H�5� *ED@A@z�%�BT��tBh��Jh���A�s�c�W�=��R�^k�������=�,��jG�Sen��S �ۻ,�K��3�N��|N�!|,�|$�ΜcB�褎wI�7�i�$E/(	��q���������U/����l��mM�˕i���r�)�H!����]ߡ,�-R�P�{�{��{��k�ec�d�4:���Z�~��?����G� �0�Re���d�
߬�SE�#��G��L�X�W��3y��Nڒ^�P&؞y��/D�L]W��ȣn�>H֦���aF񎩯/qB�	h�:�?K���U�O�g���.�nkH�����³�;*�2�3��a�!��G�`8e�5�)�-��q�������u#
��I��`�y�:����t�)Q!��S��N���k�5Ғ=Y]%>r�F����=�q�\��l��h Z����% ��@�I�]���!����	��"���!�6�@ڵ��@w���7�_�C:�M�&��-KFPf�1��!�n� =�A�ۋ�ҋ��Wyy��ӛ�p����5��I��8 ����!�D�����[Op������\���S��P��@���k_zE��I�n~�1]��lI*L~� ���R������BZ�x���p��>v�&�����ʒ���R��K��-�~�D�b�� '�<9��?��E��:'�o�����}��H�N�C�>}{J�F�iL��9��  p�Z�G���^m�J6�ӏ�e����؊�zb�4_�2������G*�.s�����}��0إ@�$��;����*ʎ<&d�g����[Q �lK��'^b�Wb�h�n0]�<�����e4���O{�:�^���I�J��5X�M@�GV��}��G��c����Z�����ѝ�N��BZ����B�	�|�R(q+z+��F+}ނ�M�jaQ�d��U�|^��g?���6��z��Y���מ�M��<�� 1h[��xu����e`����)BH�$��٘F�r1n���)/�=�qu%XC�+^2߭�R��v3K�1Cu>�=��J;Mͻ��Q����ܹ=��)Q�\�!v���SE�ξ#�gs����R�T�k��}-�i�3_�n7��)T��B�2���=N�뒼���Pza]v�m��ۛx%������/�o_�Rpd��X�ʞs{��@B��ok���N�:�J�}����Cx&�|��5J�qN�) 4�P�W�����[@��(�>WD(jd��.�)t$���Y��T��3�)%|��b������
�>MFq�=U�>~wŤ���1�\AZ(B���_�O
��x����ܰ�i�WPT��n�s�ܴ��#n�Q����!�n��۩xܔ�%�gT��Ǘ��s���H-ҫ�Tgʲ>.O����Q�a���VC=x�{�T�5�jc\��ٍ��X�-
��-[N�6x�ΕbeHvs����A��8-���	e�k����f	����\cD���P�*�:�=.fT�޺k!m�
�F��-l}�W��~��	���Y��#[�ߏ<b���ŉ/	�Emmԛ��&���ў��eԨ|��)�r�_�A��b�a�-RSkH(�	�GB�cas1�A;���U~�0���utr?�\^lK'�`C��wi�\�&���{�dAc��*S?�9����f�w��,J����^>:��,l!�8yC��<w=������))3zњ��:�l�s��:0��ycm��cB�5|����<���7k���b�ל؂�.RK}�?}�]V�����kr�����9��}���d�TT0\��x5�k�g��c2I�ӽۋKK��gU?������\Ն������*�Ŏ^��r$�zq
7vt�UyoF#�RR�wM����I����{��A�C���h��a�J�[��":e�����=8���T���?8��2%���������'r�ˋf�BZ3��BZY�h}�|
��&8�>S�.�o�ͻ���O��'������m}5�c�;X3���m�zb��9J��2R��o�����|% d�xq���_^��y������{��^�'ĿxBxI�⛇2���H�L/>���#y�����jh�~���%�z�i��$�j+�'�פi��c����N�io2j��yCM�y�)&A��|�U���U�~RH�cF�����=$U��A�����$	�����!�ǏWu5�_D�{��F��Ab�8�t����1�1�]�������s�2N����J&�B����'��4-e�*~~�וh4dF�k8SV�֖.oe��~$���v$T��O�/�R��뵠��gМ�:t�JE�Kŏ�c=�&E��i�LaZJJ�������~~Mj�"Y�)Bʱk#%�D$�?+���PX	"I���O��L���&��&�˙6V���1�k���_RR������������G?����=9�cb���ϰ�������y`���ڴL�~�q���}��Xf\mԸ�Sk�����  ���`z積1�=i��^��,,}�Si\�OĬ%RhR�t0�������w$���6J��PEͧ����'����V������X�ii���҇z�'��nP\����*�����3�����Cf�����9�S����k�����;݂�P-���4��O�'8R���Ƿtgc��ua~s�zo�^�ώ���djr%���au�gm�O�jZx`�^�˼����^��n�TD%Eȱp����g��(ی	+/���܄�h�m}��<�J�K����0�d�{L^vo��|؃�6d6�F��ϣ�����N=��ᾒ�;�F�$'����*�ǹ�a�G�5*
� �&�^i�Y���;9�>����4� �t������U	�G���/J��P���b�?��΍'�^�lPT���xM'{�?�ka����%�{.S�'[E��Z��ۛ�cy+L��ʵ�2��y�Q��ڇI�ݶzm���B��Q�Mo�X��՞�Rl����%竤b��;����0�%���	���;�̝�Ȗ~�e&���/���L|�^h'��ш�q�y�3|�1�  iX�z��\; L1 �e�̩ķ���71��qx��C&��_�,��wML����'���k?��ܨ�zb��J�C�p�C�|��#��>�8o�l�d��P�YF��wMsҞ=��h4!є�bY��棯�^X2�'m���a��dK�n�NJկO��t��ĝ�QKL��t���+��#�����"�7��\�L��%�� ��J=d��	�޽�@����Dp��14��B�>����_"�DMnWҋ�*���@���k��N&#�ʈ[�ѿxp>]��f2�)���DY}e�3��2)zQ��x"Ϟ����&@>խ^*�]L�TPX�ſ���~�w��łR�Wo���'�v�%�=�)b�׬ H���8����Q��j�"�;
�a]���nP\bb�EL��:WȲ\6Xy�f�T�"c���{�/
���������g�=b-YZ��ؓUX.��>��T��U:!��x�f9���DHL��6��)����Ʈ�:"����F.%jp�IG�d��R�&����a\z%�~e�u-�!����)�7�Xa�JGW$����e�P��&�FGǎ^��,+�R*$��Fo� �~�	f��J���<~�M�vd{E�իW�7���Ĝ�솬w���D\�1$T�	�L?~��)J�F{�1~��O�Z+T��j&�@yR��ro�G��臥�J�d
�j�ڗ��L�NTք���0 |�Z��H>���=P�"-����\*�U�k����;����N*6�P]d��ؙ�c�Qd�`�9;� �[�Q�֐u��S��O;%N�5�B�+[��Qʤ�� ��}\�yU�����s����Z�ms���cx���"g��3
O��t8'����@x���
y5��v��g2��Z��s�A�+z=��`�6�Jۮ(������I~��%H����>�/u(��Ih��ܴ)���>E���r��7�f�7�M4��3D4%�����5���)錬�L��?*���u-��q�"/�oF�v�<ο���\���Ԩ{8�E�����)&��*K;�����@�l�)���_�6��܌p?���.�H��0�}o_�'�������Pɋ�����j}$,ژ��_����n���G.Zݽ�&�s^X�ouР��855U9jy~=�F�yV�b��z��տ���zl�a����1k�[��k�ɩq\��U��߼�R�9?��df%�����5��uf�իWB�➞�x���#<k8���8e%%=�0����p4Z�:�B{�5?l���$'�[�&j��;��!i?��^���H$M��p	����A*T�â҈Q�mT�z|��GpW��L%����N�y'��͚'Tu���oJo��)�=:�C���Lׇ���M���,>4����~!����٨r@�@����|��}��?3=r�����/�����dYe�|�ʓ��C�O��	��������Ǡ����6�vj��㗷�5�{��Ւ؋�I-#L2A�ɡyMPr�gFщ��Pr���ʶ�ӂ�d��������?�N�!W��""��x�O �^&���|�v�J<�u�l�r��F9C��#����g|�M�۵�#�:��M����/���|d�����LÌ�|o�krW�w���z��>�:\����Nx;�TV�8�@<~�,�y|o?v�GF��������U����'�ċ]�Q���>3� 3���7�@�o��̟���D��Eb��ŕ7g��>D���@@P��X����E��`�V����ʛ6������63����C�7�cf@C�jt2՝#p��X ��x7ٳ~c7��1��W?��r16ˆ���3o�?�m�ZKL��*�����U��{ITm1b+����k���]|���Sp�� ��~�9�ؾ\�׌g0�������;�%����	g�UE��f�X��7��}�k`8��z%��ǧ�����r�rm���ݹ�oy��/�V+8�G�F}-7�0��~�;� ߯�V|a��4�+�z����X��M�'�c d|��[8�M�/��2�� Zெ���RN���Cq�!�/�<=Q4���.d�qOqv��+�>�_���>��R>�D~�$���1�GE,h��MP�����O��wl1���Z�3�i�� � f������V����y�?z�Z�U��\h��т�r�f7e�������u���q�[�5���O	W^^��a-�X�V�A*?�^q$.&F�3n�Vl-����d���#Q6�N��1�he�g�7�ǅQO�q���NЀ8��Y�;���69�n��z�ZQ>���!́G:^/���5�J�~nz��H|f3�mw޴��dSP|zc���KZ��m/����V����C��Z��A�b@@3	e���7"NɎ�J�˅��5�:�f_��߹Ɲ��5�w|��Jf�bW'Y�9ب�'�εz'����PΏ�z�d��74YM�*�:�܋�GG��"��+��mx2{��P�\̤�&H�4�"KS=�Ye�;�CIE6��ƴ���ҵ(D��C��H��JM+�e��:��+xݦX��9OL����"-f��@gBO?P�$����o0��"���������u���-)��wPi�ym�OТ���E%�Oa�p`A8>��	A�	~��7��P(�N�W�A�z�71�=��`6X�w2�f�BO��*	���Ϩֻ���]y#%.� ���VH�g��>,�|,V�uU� �[���P�_�eL�_��Cv^�h>�&z+��C#o)&�\[:o�3�6յ[XR����7:�5�=�ES��'�?[��`�Y���ܻ/����������g6 �52zL���^[��i�SW _�ݞ�O<���32?�8�p�&��D�&�щ�|j�scrv{@������QL���y�@Cu��G����ϿJ�/���o�)o�Y����>r����d���9�1�>�v��� j�����'�1�I��B3��Z;�?��@���m\�>����~J���%S1$���H3O���Z���#r�j��5*
��� w����V�.@�m����HVO����s�'�x��y{���=^r��Gj�U�G�"��}��Vv_I
�B��T�iv�����V�kQ��l�?E��i�[��QM0"�����1��̬�{3ѧ�\OaI�dl�$J�0��k���'B�a�' 4��))�)���]�X�)��w�߲��ON�|�@��?��Ly8C$IM�T�c1x|�3 �K5Q/[��N�����{��<v�%�uq�]]�o�܀���++�q�~$\~#!)����cO���홠�m)ҧҝWؿf�"B��6k��P��րχ�1��Wi͟�o]����-� ^ׂ=HT�2���^Ȗ�U������˼��ݰ�-.|l�=/�(59z�oJ���pY�ބ��������o]�(ص'3��ֺ����}�IB�RJ�Ѣ���52`zhH�TL�H��~�A�d��4�+t��+ی	XմT���B���[��\���cn�+u��mqwW��R���.��M�zg��4� �E��'�����l��Mtm~P�G�+����v���L��=�a}[����	SN���c�/��#�ӊ�y9����[-^�'�B�c�rNVc����xM[��%��!���.�7��3S���ӥtr	�����&#��=>VK\%���T����ƞ�w���W핖�E���P`�zHUȗ��!qK�C�(f7�Х߮+���9�a{?�B.��Т�@ѐ����U�2����uv*n�T���gJ��)��,�Σ�3,׸�2��;�ds�V�_>����`J�������w�7�j�e���>,�z�����+���N��4�(�z��I]f�S ������r�ʽ	쉶�i��]�i�댲�����rϙo�=�m�e�&#h���|�|�$�B}u&K�� ��٧B�뽖��'9u���ڕ#��s��r���]ɓ�����>"j�NQQS���Ŗ'K�V澷���tI�kv|�(>C������%$'��Sꞡ����J󐇛�z�N�	Ʊ�<K�ڼs����3N�'v������ַ����^�Y i�����H�`�����G�b�k:�:��}����\�"@�]�z�iM1�mH4��3�!��,k�Ԉ����b�_ִ��+�<7?�XCtޤ�ω0�5.��l"x�F��C�C���Lm�X̢���2w�8���i��^��>֬a6z-b�R8��d�gZ��Z��z���Q�jH��5���v8镳2ښj��֋RR�M����ץ��J�yp¶�{֮�^�b �.���7 ���O=�t����D��F��5b0G�$���y|�ܠ.-��U}����Y�[¨G��Y�bHz��K��f?M5�Y\��K��f'�������j�q p��C��H��v��K��j�6�Q��C�f��qP��Sm�d,�.�:ʘXs�F ���;�ؒ��ҽt��L�����)�M���6[��h�ëۿ���,\��c_��l.<�?�N�<��̃Tb�1�ǒ����ɂ�q1/���J䱇��tͻ�{�>c��Xr�X$˝ӌo7/on	�7[�� ߫����x��8�@��ZѷOƸ'�l7��`vR��G�P�5@f@��2�D�'6��X0�m�"O���R=Ǿe��R>:i�5�|\�r�%C���LY���y����m�-S[�V^e�*s-���_�j�f�Dآ8{B�˶���T��ĪϷZZO��k����]��M��*��� �wl��nc����5�JO������$����6�(�M+z�҂V�";���Ϡ��W�p/�d�?/�R
��ʿ��^�pH��+��*���5zd6K�	��iRe8�$l�Y�pD�O��"p#�|��CA����#T��1�C�)V��(1��Z7�upߙe��Ρ
Ł��1�o�shP����p�Gkmkjzm�z�����6��V�������5��:�3��j0���G!�1�����Ă����>�����V��������BN���K�C9�F�CS��j'�YD�����=U��z�*�o��f���.�[B�9L�~�#7�#���:�ܽu��Sr)���go���w���h�v�V�)xsʿfr�P���u�#O��v��5(��G�4~[ЪK�҄�T��xu�E�wWM��|6�R fs��)"�E�c�֏���_�Y[/�4&�|)ryef�޴��L�=d�`��A��=X�b�M6�W'>�n�>j64���P��@}�L��&��!�%t���
�}�����_C�Nq��q]G�T�G���{f��l	�b"��jc�Z籟�R'6��&|���>)*�zJ=��p/Ȩ�7���fKve���L�"�r������<.�Z{��ؑ�IR���A���>l��������6�% �r'����6�F�Lw�gm��<8=SQT�ez��\���QY���u/�Y�>;^��\Y��<�Vd^������4��*@�<u�4�[��	��U�1Z�pĺ��b�N)2uXF�]3e��Hm��=(��V/�f�n-ߔ��������n��6��:�r:����]ss�ޯ�o\m�'"OM{{�U��#����~!���t��%#�>�&�涘 �"��%�ٞ�������IZW�o@�_���XԹ�x� �1	�׹�ܼ��!���N; �*��A�>�j�B�<�9zۦ����+ut�>ɘ
۽o�-��q�����*�Dŷ�b��@+��)��K��y�[�/GQ׈WRS���x#�Ej��Z��㏻�����r��]Ex"#�"*�S�N�-�Ddk��g�#j�Ï��P���s���\�-���˴'ּ��tЇk/0���6�U��eA��>�s���?�9*�ϡ���;rh�.jz�{n���,�#�|��l�c5	A�o�
������67���e������7�p�	Uz�2;��I���,Y�=\WO�YEc�ײ�ȥ�C'4��X(��f��k�dT�E)��:r�i�nX�V��^�s�Q�����Hl=q�wz=Qk�t�
�z�P>�EA���:+�U��a�о�}��ﰠ���-�@$�����\��<9��%�$�s
��+���P��,�R�ʝ2\��0�}�J�f��Ipꨣ7��x�@�؉Y�������g�o߰��ի�S��hV��Y��=bZ�{�i�t�&F�K�/�u���t�3&��\b����V���W�fN8z�$C������#~͓�\��

O�~���<E/]	DY��P�<���d8i�H�|E���m��-A6唦Ӻz�^w��y0.��@�~��5h�`�@���VՍ��/�/6R博�����y׋x��#�3 ��͌���Vz�����#�}���4;�!c�R�TD)�.����	��-aL�g�^= "�y[��I	�Ҝy(+�z����d�Cl{Ֆ�F(�/_�7;r4M���$$��3h���1��L<u˧(t�oe@��a���ٝ��MZ�F��A�
ݗ�{�R�W�X}Ƙg�j��R�u��k�1M�A�ޯ�0_?Øz!1c�V�"���v)��?z0������oЀ?l00���'R�mҔ5H[���*`�~��>lv4G�1q�7L�叙(v����3_�o���u|��?~t,ț}C_, �sG핻��g\,ʎ��s�ؗ�8��p�r��&o��2/�u��'���o�q�T:zY��f�_��c���kN�V(��ijT�5��'�"4 Q��*���\�l�B�y6�^��#EV�H¯j�����g�Y՞���U��;����\��<�����]'q����yĩ����݌gsq�(�`�J���qM�MI,�h�N�ؗnD�Y�ln^��(�i�����PBXX݃\���b9����I��ӫ|$׶K&�3�\ba����#e*��7Vk*-5m2 +��}����fc>����U*f`6Y�"����)��6�Z
툅ו��/T0�0��>G:	z7h08%�Զ�)?�r���{�S	j��LM� 4?HW���`_h�s��I@��Qs���i1sk�Y�Y&\��}���2 ��(�pRDl�܋�d��r@6E�)���7!d����r�S#x<N��.ܽJ����0٨���j�-8]mt�(�Th�Nbn������~���}vP��-����%�Y�%]�� ��tg#�ܥ�-���Q	.բi��>߫���Z�h�d� vW�y"nrʱ��g��x�ku���X��a��%��Ӄ���%�ЁXTV ƇP�U�Z���3��h��얃�����f5��	_�E�V�t2�P{�^�v)��X�?ȷ=�r
뫷[,@ Y�; �T���޴Gդ%��Ѐ�;qУ Z�+ܓ}4J6vP.;9LAS#.S%��[����ljA�j�y��q]D�)�k]U�������79����|`���J:��}n�r��.ט��[L��CĆc�Fu�;�+f���"��aX�^�� �+��̩ʻ�'�� �g�8�4f�y˶�t�?�c�|�.i��(r�
��d6Y�܂�]��S)!���[d��M����p�ʖN=K7�Y
�8W+�n��%yLz��:�ϝ�����I�(��Z�$= ��k����m�q����X�1��r��ͨ����,���q�?��ȓǜ	Ks�|� Y����8��\Ir���U��J�3$�YЬ��$����('^����o�(�K�I]����x9��-��-&�e�J��[�������J�))���Z�0�+P�}��.��f@-���Gg��"�^HdVk��Y�|X�f��$k� �i;�Mk��OGj �9��ǋ Ӌ�%|i�\�UW$�?Yt����aZ�>�4p̕x�f�asҜ+��|t|)M�[B�q���o�|�Sļ��T/2�j�\}*���`RO/J�f%1���͛@��;�8����*����Ý=��wg�u�s1����f��Aɢ�n���.�IO����@����e�i3�e�ZX�����,,����%�cҦ�<��Hhn�In�d9�6`�z#�؂%�'È�-�F�7��ʫ/:��@��q�)�8/Ib�-(��:�J��_�o����K�#�!�uJ/��A`��vvIj��S���%�+Uc~Evj��d��c��ꌵ��>�t��2�����`����<Q0����`j�{|l�����zba]�E��!�:=�νSdKy�o�/:,�Ald 9�돦ٸnG��;k�� ��l���P���t��$����y!r�KƐb�yi�5���ю"��	a0�p8�u�ԡ���p���T�0��#�'��
��<K1=9��/<MJ��/\��^ �����OYn��o�����"v���[����Y���ef�\�u�}�l�A12�i�.-�t�g#B,ފ�pOdn%�ؓ�"u?������k��a�1���B�*�+���ð���
au�Y��|��w�5Tu��T]f�}�Jº�- ��N��L���/Tz�њk�^���O�{�%e���p�S)BH;% �<ۭ`5�B�S ����Q������mx�^ǉ�����E�3���F5�*�C}r����bC"�Zs'lȁq�LC/['��?+�u�0���Xn�:?�u���զ�Y�S\N'���e�2�Yv���F��n><^}���O3�Z��]��	���+'}�G�5��{p3>�Z�&{g�Z���|���mJ��^/�p;5!�
%�}�g�`�"�7��HgkÃ�D��Zk=��Zh}��OO�˫NL|T�뿙���������8y��+��.����k����u��AK�ˮw���B�3�t�y&�����8n����ϛ�U�&�����ǢN:��%xN	�n�%Í �1VӬ\�� Q_9������U�O�m_NGӏ�[�vB��mJ�^��@Ң�K�X�1����!��O�B�S���"P4��Z�O�Vf��R��{���*����ߢф�
�==���F��&j��;7X���#3�S���UK����gS��%yf��$CѦ�7����������\ � �W����ޙ�������A���c��T��z���_�vK��]ݐ���:��n����Y�(���k����sJ�rͲ�����t��j*MJ\\��[����׸�^�.|��
��6xic�����p�#kp����][�V�H|�^��]qau��R�-��nUWO�P5o�#o�zm�.P���Y�Թgz�Ɏ�j�_a�Z1��׽����u@v�@��������H��ck��W.~;K+Y�/�l��3]jg�=�S$2�D�:��+�I'[����H��S1@�ѱ�k#�y���7A� �@kbN�6��:���ϫI�F(��{K�q�ڵ��)vI�6>�<�%�?�'=�cz��܌�p 1�<c����l�K����L�Abꑁc�'[w
��5q�D�)�E(U��像�[3p��|b&�~'�r�GQ�g�{O_4��ċ��f��P䰿IS��W��ȱ{M�Cʟ~D3K�0�)ּ{ȍ��,:�'���g�Y�rzR��ԇ�6┍8�A���z���:����mJ�&����Zʺ�B~۪���=L:<*I�z "0�"g���oO�~-ɥfw�csQ3�DhOʰ>��KGX�`��P���ZY��m>re�lÏgD4�7,����0oee�Z޹Mw�2�q�,N#4���6�3+�����O;���1(���)��~v�C�UL�Cj��gN>�ݾ��}w��)y^���QD��L��s����D�z��	�������rS|m�flC��_9�B]�+��Y���&���+r��&8��ϫ�}q�q��Ag��a��3�⛱Z(S�����r��p�9e�|M`�@;`�?����B�Dg�w.�A2�d�,'�J	�e�D*��wbT*45��z�`�C�{ WSRЉ1k�b�#��zN֨j�g�R�ȮR� X��=5�ed�;� �n�?:����=x+�AU�h���ˤ?���a6��7�*���!o�lv0�ۧ
0�)V{�xn����%���?�.xbtӛ� 
%.}sAN��k�!������p^^���Į��EYC���j���R�7Z<?��:���QK#3��-c���}Ѐ�rM%6ȑk�� 7M�����0HR�`(�[�"�#���-�Ε%5������YU�K<��n���,ֳ�|zp�\X�����6��jOj��R_�/$X� ����eA�D'//<���$��l�#��ݳ����C��A�C#D�������?�qD[�A�����xK��k��1�O�է�̲��Ջ�}އQ�e.Q:�HJ�Lx�|`������oT%{��C˴>����%���6�Ꞇ<eY/μK@����o�&ce������X��i�,	m��k��}^�h1s�K�n�>��М�I�]k>_�$���y��&Zp�;��#�v�o�+�����p��0�`�=B����������qH]RK]��_>O@]��Y�֦M�ȱEN�r<qi�:��Z i Q6��lX�%`;np(j�3�M�����/ii% ����il�Z��b9��8�f=�4hD�����<���:����Ma���!a��W��(�л��gV&NEs�ΏZg���Ż�|�˃�шj<�:�U��1I�aH�퟿,���Ԏ���"��N��w�?���\�h�y`��Lf#��m�*�Q�^��ngq8K4/��������t���;���
��X>Q��h��JZ@&�y@ܯ������ӆ@�H\\���%'6���5'������)�D$1����!�v����=�IH�D�h���҃����B��q�B;rQR�H��=c��EƤDdo�Hz�.Q����\�A��N�[{�¯i�۞�;��(���E��f}��vL�^� �0$���!�z$ �O!�Օʫ�T�,
�Y
C^��wۀ���O� ^�e�e��b��/���m���l�l��μQ�L�e��Ņ�ZS�ev��Zq=���nR���x���ݭ}�,����� '�R���CUPb�ã�X��5�ئ7���]�ρ��m#=0s���`�������������s) �o�K 2��}P���� &i:�����j�p��(�媆m��m�^���̃�O�b(OB!�3�qV�] ��.*�� :����G|n	����h�I{ɻkn(��5�mr��i�v�����W`��,��cR�>*�k�'G�ڀ{��w1�r�kʟB3�s=��*w����� d���������
�t�y;mh����d]��ٸ��������-Q�M�Q1WH	�A�x����;�#E,�eDD��5��z��rVX�������B��ܛ'�'����w��V���}*�:io#֕���Z�A&���c�LV������}������.;�/С��K�}�Tr�8�.��7��M�L��(����'�vC|��#}T%�J��9a��H�%��{忥Z�Ԉ�Ă���c��ּ�[����	�`�Õ��rb`�^�4m5���&:�^���������7?�76�%G�[�m���i\h����X/0�E�Ը��D���y̩�ܻ�J�3:�2#�> ��Y���Z���j;DW����7�q��-��N�'c]x 8
��a:X !�(K�{̀,U�K9|ZI�$��O���8)��"��0�o��po~���c>$���E�H�����-p��^w���~{A�#N����ö���󢉭&&q/�����<�Q��u����C6���*HM�:��T��]Zx�<�h>���1F��`)��T�ڋ�Y�o�^|�u�I��<��ܰ�D^d�@>����c!�ί����r���Y:��cʒ��{�˔�=D��X�������T�[}�R=�" ^���bV�Y��~Xm����RD�0G��O���ަ�9�� �i��ვ�@׉S�n<���N������҄���/�U�ИD�NiȌ�}d�Ɋ_|,��1UL��@tF;'.��_��涴��8(Vz֭׊8u�<ꨅ�댙�Xq<n��Z�[0�XX؜�c��<8��V�c���w�*�R�@���2���~" _�
l8 ���_�%h�c �Hu��K����LL��
x��L��9�>?G]�xϒ��^X�X�B��W[<yF��	��*���I�����pߡW��Q��i�@���#�h��3��~�8�����P�jP���1ſg���Ʀ�򫝾%V�G���$�-��sӬOM7�p�q�����jL��>��AY
��?��z��"H����(on��#�|'���c	3��bL|�4ڬ>?�5S�eQ4��UTT�A��~��l��w]�z��'��mʈ]#��!~p�L�a�,��+�س��kޒ����V&�ꟀGiL�*�{拈�a�?���F�l�c�2��敟J����[��>:<�iR�&�P��e����4���99����&�0��}����������t�º�����T�Uʆ�MK�${u�Ø��@`�1�{J��U�&Z��٧�-�V�.ϳ��~���A����LNJ���M�M�X�1W�V�x�����k�Ap�có"u~��u��@7�M�,������j� }������s���=�Ԣ�28�#f� ��������J�9x�@�ğ��P�[���\�3i��hqr�2��wx���l~l�*KV�{���c/��,��F_�4�\�ތ.0�,��U����8%��I6�^��U��>�|�G��r����S�l�N�x���Fh��|�1p�*��X^�s�Q񊕈�=����	����\b!c[�����{���XU��2��v[�65�Y,����z|M�у��������`��p]���p�=�\!v�7��<"�C��}�<��ܐ�v�X�:���s��;���4�33�z�Չ�_�B�����=8<�1�}����6@���Y��x� �D-K��3����ދ���˵��Q����"`������ƣ�!��LK�C���{"O�m�҇���j��	x]�~wI�F���O�|�wן]�|!����+v����$ro��5��/���]
yCr{`���Y�I��9�˳��W^����0���|��2�o9�	�����D�B���T���7��iK_�t#�Kt��1{n�-E�O�Au9h���,W7/y��'�/=�����;�֋fB��u�,Ά�v�8��0Jy�T��ޅx|������'�q���r�IM����������*��t����}C	��I�H��[�~?���3њ��Q�Y�'�<��� �v�:go��W+��V�¸�<[JyZϥ���_Y�H�m�|fq9�b�0]�9Cȗ@�rUk��wi��U��SPý�����'�蛥=�;�B�		��x(��}	)�W���u��]�F��Y�k4���V|fu�}|5�ה�y3�sk�B������ ����0>���Ծ�v"a�󷫼��.-����f�]�u�C�����?�tS�
_����[�Y/G&�Yq����cPa�TA2�Ǫ�����ڕ��?�|���jT���.p�0弛5�P���q�9�[o�N̟��(Έ����~����=��3^���ꭙ�.�АKb"�T���a��w�����Ņ%;�\�LYB��"L�i��L潧Z�o�2o��8��|�*�ǁ�����n{d��&����}VV"����*�"j���+�����>�$XZV��s�?�96>��ߗ�2Um��]�:�,�%����������z�����c�/"*����+�:��(�� ���w柽�����y�tu��%��������v�����
�X���tp�[�'����7������n��:�PO���}+������x����Ľ�2��>�ۖ�ou!c�v�����{�!|�������M6�q�������Tj�Ԥg�Gm�������j�އ������CBZB��������K����n�z������l�>g�Z�z�}�g7Hg.��ұi�ӐHd���م}���=c�ՋE~�),ȫ]�-�W�u�NN��u��"8�h
��y}@���G�������X����IXO��JSF \�8�o��Jr,���O����0��U(�@��y��^s�T.�s�n��/S1�Svھ,gsqÛ�y{6��� ;�r���������c������X3�9��s��'�p�1p����36:��9:�F~n�jd���*�qWo&��nWp��]��S�+3��L��	�=|��]�>�-��M��]o�~Y�U�\2��)G����"��`���d��=�`oc����+Wc��O`|�<o��U'�!�� ��c}a��\�(��,3�g+h=���ɨ�L�I�w���(�k2�A��(b�FEj"�&T݌����c���F�ᱣ�cC��+K��4#�� b0nK#65���Ǝ����z���Ȟ�0����o^5獽C#,�¶�bP?	�j�R6����Ց�s�ҟ��4ᒐ�D��CJ*Xo�k����%�<$��Ƹ��+��(O�s�j6$�U�F>��.A�\s{�7%��yy�(�)l�=�B�=���=���y{�e-AxrG0�Q�����k�*��a^�]��f{��砗�ܪ~H_j�l����lg%7��oʠN�����]��~�zywhs�*F7�:��wh�����d� �ϥp���Dk�5w�I���N��N��N`�\�n/�,�-V�P��6�42���&���o;�	�GY��t;�y8#K�8�	�a���.��&ێ�_��<�ir�׊]��;��\!3��z�l���ptG��)rI��֢A
�
~g��VBn�B�F:�L?�/93�$;�����dN���@ܿ'G�5��7c�=Mln��g�Gw��Ǽ�����M^����S���ɴ$�+i<.x�C��u{��:p6� BC]��LBFBY���pa����y{ȅԿM�]5����[Ն�M�������4�#g���X�U�fg-ߞjܞ�8[/�A��D�樉�$l�̐ۈ�m���r�~�����������6�nd�/u�z��߫Ȍ��6?�
A�['4��D'���e\�l�:`��܂�����Dl����|~p������D��[�l퀻rff]�ן
l-���s�`*�����uM���2��I'��$R	C`��d������֣7�_*`@�6GQ�e�!i4'_6��(d�֓96��;H���S��N.] $�	2'�@��4�18O�W�n��T�	0}XNB0_��@��]0�Id�n�`-�o0�`Q���+��J��U<<<��)H�Ŕ�uY[��fw�}��������R�Ep�D��).��}���,+)=D ��v>�b
m,�p�'kp&h�-�4�0G����S�hmW����>��]U�wb�eb�����K�Vפ���{��Z��ͼC^�H��"i�}�$�;t[Zc�u���<˨���ͣ�Tkzkw���'�{!D�-�ďS�ꪂ9��D{t����o�9�̊IΤ���[Xj��Nv�d����x�۷�]�ɷ�	L��K��GX߶�¢��r�M
��[@tM�,"�-��a۵?�!�R��Hd�yو�:WO��8[��0�/S���ъ�,�dE��T�*���YBrYllB�h�./o���Kt���ۣ�-���T9x���'~��i��:e�K,� `�0��0�tȞ7=��m�vo~����O��,쁙QUkc&�S��E��������=YHR�
���g�n�lgoP�w�[�@�ɲ�B�������Ê�%�(��6��=�k��jg�V�l��K����JY�H�{�pp���C���2�"m��a�?w>i�xq��D� �u�'UB���ձ�L)�|�W�Qgs+��+Ԛ�L7M�ə�yD��,��/-�fy��O�|��d5#[3h�D:��U������	��+m�@,(�ѫ�?q�O��y���E�30/ �������BWS�Kq�#�07fhfUQ[Aǟ빧��7Z=��Y~U����IԷgaA�x��w�9=���-��w���FD ·2��4��so����)B5�R����	�'�cӉk����3�<p-��|k�=_x#�Վ��7��Tٳ����j����o�ShT���@_$B���|�06&����Y���#���>	�t���0���n��>���O�6�Wa�0�-T<
�(��}gg�ӵ�C������H�%|��j�ɿW�P{���N��o�ה�<�;��u�}_�j�]]���{�:��l��ν���F�׮�ec>���mӢ�O"gy5K>�}�`�|L��	��0�s^q����^^K��LY����Zyj�]|�O�^�w��v1q��'k���y�Qo�v�s�n+K��МI� �DQugd�F�����"��oBh�9�M���UR;�j2.kԷ8E�;p#ր]�.T�j0��E ���}Y��'[�Q��P���A?�G%P���c!�{`�nwP��1�&���{t׈����)��E�/O^֏`�?&�>7M�ea�y���J?6\��[�e�2�,�H ��5�;]�����/_6�,��ڮ)J}���*'6��س���N>�����0%Lz4ʙW�O�ȵ�>��v��d�@?B"����4�|�uӏk���6�b�hw�$[@�y�}�g7M}v�,V�����tQNd��?�!�ct5�w'��ZX4�4On�45��ka���@�Z�#γü�á�~���Ey4҅a,Zn�xQ�6.WA��?��L�
�d�A$Ғhv�� �uO�3y��9���L����_��Ĳ��F����=��ҧg&-�03����K�ӎ��| +Jq)ۨ��
X�u����Ϟu�hV]���ă������1\�Wl��@�!v�)m���B�J) "vMu#Xq?����l�fFZT�;����)B�"�����)}$i!�!Ao �����7�l�R;�k6[ݠy�Y�8��VEV^z��i�����7�U�@L�ټ�� W��.p�:���p���J��K����]|�P
~��N;(x `�1�ۊ������6b�;;��S�Mr���N�p}b�%N	�M��	��	�&��b���78��n0��=�;i��"u.�����e� '�[lR�D�R�a�F�zr��9p�����ד��U?K����>��v�:,���B���{b@��m��,�?Z�\Sߑ52C���� �ʼAc�8�F8i{|�X�$�U��d�*Rx�\�cY�z˅�ADozcǼ~;{"j��Ʌ\�8s�����7�K_3�m�q�b ��syXOl��
��!t����`�����#ܚ�/:�~s�^�����6�������wM}�W���+�L�_ฟ�DK��I�ڝ�2�ǃ�nb�2��P�����嘆'�_8�~���*�G͆�FYȸr��Z���p׳ċ����٭��C�8�?�2D>ڷ��]i��V7�������U`*�Ɖ�b=�->X<c�ւ�ر����p%���ʷ�kPW��\���1v$)���wj���G�����yu��ـ\BЕS�(UM����b�Xzz�7Ooiؽ��!$_�n��@.�"�X�\x8|P�:^$H�Z�����w��� �;���
���\���R%CZ�`X��-�~��{eu1�F}�H/1��z&%G���uh�����b,ZF%�`�Ob<E�/�e=�J�����������Nͫ�;߂��ƞ��+�߃sUԽ��K��1e�v�����"A��D��L	���(�j*P�T���m��d��P�}r�YFY�#D��~\��)I�tFU��slF#�`��m�h�Hx�^�(ke_�"��g��o�WVĽ^.��0�"9��7� �-�H�Y���$�*â���{.(�M6��gv��2t_�3?'����DG@��ڸ�j���Ȕ�m���S�y�Y�O�շ1�D�ٸ�A\m�>�K=�� �/s�r�����/��j$ow��:���0��-
�,6�&I�+ �-ߦ��уԮ�? m
~�F'��� ��i�Di���Ĭk~�{�7��O��/� _��-��;��z)�fu�	����H;�9,��	�{����Y��.�����! +&�f#ؕ�����9�Z~�����2Hfd��_��L瞂�
k߀��(-�5��B����]ٗ^������$��n.���W����H�<�������?3/k?`	h�L�����Pey]�UN���N� ��vGO�c�p{��@^\gȻ���&�oU9ʮH>NIj���`"����j��΄��	kňj��ͲǼ�S��$� ��q���*T��oŶ�ZT�@e����S�蔄�cPh����vnET���J����9���VX�M��[�J/:�ՠ�J�w���!=���#*Z����ץ�.];Olf�7�!�l-�pC� Ġ\��C$���m��g�c���c�7K'ֺ��R=F)�PN����:}���O�,a�TvW�UN~�%�F�����{�p��:�My$�FI)f��p��w�-$!����ɧ}��̊�à���(���E�AF���N�ICc�3|��"-;4fC�G�a���s$�㺳�s3�|ͯxݶ�u[�A��܏���sւ��z�'��c�Ľ�]�d"�m�.�IRS��]����C���������^�.Wն�2)7�yp�L_c��A��_��ԇ���G��PB�?��پ�#��s�9�^���[͇U�6~�m�R'B	hJ|~0I��
{� 5�k�h���"��C�#拧'
>i~L�
��z�>ilM�?��+���I���h?�!���7S����R�6�'nK>4�IF/I�gݹfl%`:�f�T<�W��.�q�::r��"ϛ����PU~���P�W����9��3Ő���f7\U}��h&�x�S����N����v
�y��;�g^۠�,yl��`���ʸv�dK�s;�h���������K�Z�#_�=���I��|Ƅ�N�1�|uC�L�5��ҀH�@5"F�H��DZ�{���9��h��,V,�}]E�y:E��������7�y�'�WB������OZ2���˲3R��B�/o��W��|jǝ6�1��<Y5��.����m���P5Xt�����p/�{�d��TWs~[c3�I�"�lUM�����Y�B�99� �'�[������V:�q�`�\���08�A��Lr1 ���R��{���ueTٮd��a��w�Q�{�<�a�0�zq6�R���ն�=��֊��PM+,��&QE)A��L���][l7g^�4�O�qC�ダ���*�ߥ�������n�V��A���Ő��ެ/�5D|a�_����L��8�m��$�x�d;�yh�]W�t��r�<A;��ߺ�ʧ"M����p��&W�݊����_
 ���G����a2�f(��-�2�z��t�f�.�_���r�4p��u4�/$Fo`z�S�U@��B���U�&ig�y4 P�n�_�u�Qc�W=n/9�h;�6��Ah��X1Ga��M��]�����^�)��kWH�Rl23YI�]��_�)�q�A�-�3��n4W�	O����z'}ї���FV@�]�F��1�Ms+ �<�����y���E.�&s�{�b4���p����x�����n��ǰ��A���5��oY�@�O�/-[vP�tҧZEt~�-F�3�Yz���@����_݊֩���Nt8rK���s-92)j��.�������%���<4����j)7B�k�\w�o�y)EQ�S��o/b�4����fYT��k��E:�IY58\�����|Jn����`M�G�������2�(Mb�ț�G|���F0�ϳX)u��_���
��;�;:�oN��|N�R�6K����w�ܤ���=V ��s"#S���hm?�~�B�c���s-�M
�0X�A	Y�F�#�6�I�T^s~��N���$�}� ��e�Q�%
�߈���}
���0&]l��_��o�ѯ��1�* �1b�X��u%ō���90���?Rwf#)��S%ʔFbڡ'�Fm~�==fb�0��PMᯡ�'㷹��H��F�IE�탓|�fw�[�>X�[ۼK&��`�
Y������۵y���
SMq��v��eo]��=qPw�{��Ğ<>.��/
Rf�v��vms�����*�%ƥF|el0\_�X+��-��Z����:꥝�˸�E���f˾@�7�%ˬ������h
F�U�D��\��^����l�`Q�l���%u���lAۦ��F����}�>��~�;KL8������ oto�*}��-���@��A�vm��m���}玏���w���n�K��)	x/Pëg�u�q������hB�����b��w��*y�\�ٟ��)(3!չfSƄ�u:�j"�� h�?��W(x�|uz���w����C'�)B�``oݺWc��X���߳��<���������P�
���=��/_~���F�]�[�CiV[j/��u\�{��3X�bd��.cP�R3bM��V��K�6�l&�>W.�a���wj�1�ֲ�����LP���f�vt��{(���aHr(_��Z,�9'E؝j̀��і~k��t�+�89��*Z֙~� ��͌@��Xo0��E��X_�������D'ڼ9��c�
C���ˮ��M�ޫr� �C'y�M�1����i������f�	�����7&0��{p3�L�)5a�wu�g����3H	�!��?gҘ(�q`�R�ɇ�5�27|���)Z��P�bp�&4'�V����C�x�/�5��lX��gS�`W���Lz��
6��bQ �4�z�T�����@,��TLg����[�z�PD��%D�%f����ڵ瘀n0\+g��<c�l�������%�7�~N��A(351d���.���)Ӂl��DaA�/����Oy�2��1ƾ,i��2*�s�W.KW;%3x���0ơҽ���A�%�O���TdG6Xs��X�H�,,���ڂh���v+�!��l��e&�%X��~�_��� ������>�5���om����n�%4Ja�P���R##d�6�jG�"*�$��q��?�~F�a�=��wB��X����GK�(������j{��e+�:��xV$��i��R_���w�]2 ;�d����;d���\���[�]�u#.�m����>��ʇ�I�PQ���5{�[T���=i^�KٕP��W*@c�:���mU]6�}�ۮc�i!�W!��lB��C�3=������ǒ��O%�����m�vL�ؑlWG����7S��^����3����)|�Yh9�c��$���[�&P-�u;ݺ�7�R.��E9�@N�� ��L̃3ϧKU�:�����3���N�a5�'�"(�e����OL�����H:>Ó~��[[��f�Uٷ��7��H�Ѐ�G�<���▙�Q6u����p��2�'u8��1�;�����f��e;��p٧$7�hv(ӈ�X��^1��?��:-,��"*U���Y�u�ܐ���fm�Et���}@�T�U	��|*~Y�A$,s����lGf��t�j�u�~��\I���Kt��-En�:�'��\�����c����m��J��ã���wM�u>�]�2(J���䜷��4)�u?���EZW3�]���W������_t���eQT����������}���c��ټ�uؾ×w?��#��j��;<\��({����l|]�����/��a�*w�^�ႇW`�H{�1�4_��0 b	�?V���I��#O�u���}��F7��^ui�����
8�T������hIy��Ke�mQt�_/P1���Q�;���j���K����}�n��X cCㄮ;�(��)D��cSr���%r�)�	S��S*Q�mMd<�����׹q8���q�r�6xx�]��z�A�����7���8
Z�������[k(��_��W�k~b�f��+�,>�2�hWU��_h������E'u���Ht��u�2����7n����y�Hf����Hbݶ_#�F0�o~�}��i'���~`Ct@[�Y<R}���o��u�����2��	o��䩔���+�qjޮ���X��๶9CjLk�3v$��L�s���fWYy��<M�oT��n�I�6V���m�nş�	qMvS(��g{.P�/��Q���?��#�%zN�K�����!y=K��q>��1�<���}:}QR��X����ѷ�����I`b�_�"h�"MW�JX�8#fd&�o[�M'L�bR>��EQr��w�B�,��r3ʁ��ugv��^�)��:�b|ڗ�Z��'�@�1t#;aF���ê`^��P�D�����8�l�2�]HqWa�ňQ��h*�� Wzm<��<yd�
���S9XKɕ^P � ������C�Q�����`4[0 e�o�hj�n9R������v�Q�"���8��}�auT=;wd�_@GM~��W�3���^����<�}G�%�מ��YO;V)Nj� �����AqPڥ��^�%��9�3.)3`MH�������A�r_(Ťy��-c����������K��bN��� ��� �Ή�XG����g�垉��=IJ�:�D��r�� #���1����<<�������2 B��_D�9y��+x��CG�9���X���͝ɲ�<���_���ۻ�C>sb�P�9�bp��j�'f��Q����Ic^�z�����{0��Χ8�fU��҄7ߧُ^.�~p��\=�~�3�O)t|$��FMDfV�!yn�M_��P��C�'���w�x���u�k����(ll:�@^o�z���O��6Ul���)�g��W׺d��h@\�"�@��@d�{F�\�~�h�z�`��(8����@n�~�Q���M����G�q�\�JBr���C���~*�?+�� �uW��g~p�&�sh��_Z,�`������K�W�h��C�՜�|��;��ěg܁+��jQEU��r�Y������^j�<>�2���݈��~h
I�V&� "SRE�g�%��Gm���a���Q~�0���+�!�����K� y艡�$�YG3�P�{��>tdGSC�p�;)7�;iGE������5{50�@��7��hG�_����{���!������1W��w���>�|н�&RWJd	eJM���d�?��K T9'Ņ���-�O�*x� <�-ҽ�+"��s�A.q{��r�{M�-P�	�O�y0�I�u���i�=IL�}v򢎲���	���Ɨ/�P�!�@!�?[�M㹙l#}>�`U�~�$�Lqw�G�IS��] �Spg)���A�c۴��p�@$xB�����ht1U��:@�����#�*����g��y���k�DB�+�l�kx
C�T>cqܰ�Sd��:�eB�v�i���Ƙ���O�ȟM����3��ڷ�!���J�q-&[�[��Г9��TE���i��* ���D�{T���ն#�ҕ[�@<���n�*�8��s�m�����B�2�pD�S��C�lf��a9�,�P}���C�0(E��:��ˌ���C���5��Fe����&�_z�R�e#�%�I�ք*�v�+$�S�7e��ۘgs�[lvsD�i\��6���{OO���5�\!@�Q�T-��<�7-*��n�<<���Ud�g�����)̀�V�,�P��|{>�I�f)�(��ϟK;������B��<}�1<�9���D<|�0�ؔ�'�&�1��0^(��?��.Q3��˩ӂx��=zh�2���4?&��aL��P�?�PQ��o��`�l�L���D�A �[�=D ,K�,��Ds���>@�ޣ�`R�����8Ƚ���t�=;����\�R 	�"�F���EA����<�zLY��G!#a\��
O���j�=�Ӻ~���k��~�ШΘ[a���z�OU-�jY�;${y�ѥ��1--��'_��X2)>9),�k�%�f��毷����]X�𱤫\��y�x!z��l��
��b&�y�e���L8�l�Z4f���3�D�M� �E�҉��Y(�\"ͳOz��#��ۄxԻ�����Ӵ��C���,M���<UX5�%O�ڈ�lo��UU��%
T���7��������_�y�yPZ��$����o&�WvN�%�Q/�`��O
�����U����x�S}0�so�&8 n�R؛G��mz�oOSyND�7�|�a�4ko��`�����)R�ǰIˑH3=�p����R�����ת�xmm��� -Y����� P��>`�0q��0ڒ��xo;�V���զ;�i'Pg����ÈG���[1Fw��b������%���/��!O�q�*�o���u�
��+�$�F��tH�گ 1��X������?_T�'��`eR(�ebSq�g�Z�nF�y%邾�����C&x���kU�����ܣHM���9B���i��*.�*K��s�dЖ�\q�ڍL��W�����xa�w����L�����̯��R����N��������5��s�I�X!t��fU��2@�Cm��sN�џ��X��x�*KO�3� ��Vi9N��� X��BOa!>j|c"�}&��if����5b�C6��j�ɑ���=%q1#6�˲�Ȉ�S2M5��H��8���	��?�AD���u���'�,t�&��`Y����}�:���R �W������q�<�eeG���R3�����l:���$��$ٟJ0`'�����	&�0=�ⳋ4{�@�d����&�u���.�-�/Gz��K#.�rh��",��'��Roa��?�0`+x�@�w��&��r����;D�h7�Ę�����{�I�����k��Vb����%�ט[M��7$�k7\�����A�	h ��D��F��.b�#�gu@��Gx�<PC{>uxK\�-ፎ�*�k���;އ���]+0��^��8��,�`;X�qi\��/�Q�̶
aRa�X����㍆47�Ym*��H�KW,O�zY��4�˜�H��^g���A��<��)�����J*�Vs�}:t�т὘��e���L1I�D�1y>ܤGK�V���ϩ�2�OCP��2��y��h4�1��J	qīCf��D�Fv���`�a��	pX�} �U�q!�����LZB"�$�f��?��<�8k-9���S��9GҪ�Ԝ7̠��C��p��.���6Г������=�>�p��RQ��7�g�e�:?���|"w2��h&m<3`z�q���:�B��(��c|�w�Qu~R���F�7�L�[6�C�`���<~�0f�W�#h�iy��%<2�9��L-6�u��F�pa�h����M�] ֪������i��T� �z�� ���B�coV��Z���[U�k\ub��/�HrA�ӡ){QSt��ZfP<����T��1�{�����`�/5K�<�G��"�]����,��s�c8�'�\N�pRu-�x�6�����Cc�O(�e��/ŏ8��ZD��V_ߑUD�2��E���".���$N�A�t�j�)Y �_���՝/�&�+����S	٢����g�TE`Hv's�w�c��@���K.� �M�9�Z�T	�(��g�Re������!����6
�?+'g\�d�G�par�y��T�Uz���ɚ\�T��l�Hh�h�}0�쥝��ěol��+�v}�-��rz��6={顗ƈ�+���R���!����+��}u"+�Z4�<+SV���ό��7��eI��߮hg5{ϞJ���	ZҰ�跪Ȥ�� �ݡ7����;�-��?+jɌ;�������	'\8�Y�����5%��7o�.t�~2Mp�a��mB������nd
�F����c		\|]�y�jn��&}(�6�~���O�9�H ,����5V	b/q����$��9Č'���(9�E-�;3�+n¢J4��2�q[���&�#�YˌS�/_*��Y�aø�s�����i�[rF5�[[9L����@<�y��VZ6Z(P�M|)��L��*g7�2�2�WD��̐���8����Y���#����+��M.|��+�Ay���;����X�faE�o'^=�S��(�$�Z����B���>Ξ9��v����Ih����f�w�rS�3��[�2��` UUǢ>��GB\�m�zx����L�7l@f9��"M��_=�
hv�1Lr[��6  xt���7C��^݈�\b� E�Aj�4��ʨsy����.�S�z�8��oZ��Q����������#O����a}��~�o!����׺5$��Gb�K�����hk!���]�������� I���:��H�W�B��K^����>�eO����?�DKI��y�?I�m��x��� g�@'}I�	l����闁�H{�9�[^�<��V�5�c�C�T�����5/�Xi�3c�WU>�~��u�����[�����IE��I73��ZS�G�w/�+�i�y��u�p�"�E�N56�2��#�}�4 ��-�J��Ɵ~	{;��^>��X�?@��!_���|��@��B4�w�-�'�cm���B���+��HI��wD5:�.��
���7I�!Ϊ!N�Xԫ3�t��Xf�͖}�d��Xz��KHX��|Oˬ�� ��D	AHz������t?θ�ߣ�>h�\��A��<a'C(<A:ݏ����'	��	aj=���Q�N�~y�|`��'�-ޢ	��5�^���6�@���&U�ϕ]��JG�O<ѶwV��L�$8�����Q�ڂ������`g� '}	����̃krI}yH���i�Q�C�g\��27؏;ռ,�{oY �P/�������$���Q��1O�M*�*fi��7I_���Š�1(� g���-�!�;��ǻ7K���~��6�������|�c����m��B�� '
�~n��X��O����w��H��;�9 �'+�=>�y�+�'�d��0��`\�U�3���>v��#�õ�|��3f&��~��	�6��t����(����rT]Y����Q���O�ʁ1p�Z,�r8��t?ٸ��*A�D�G��/���S��!N��W��y����Z�����|̝���,i�x��W�a��h2��4=��߿?��ś���`0!����]�9;!�-���iC�J,M�MY�}����a�gk20C�������:���: �RvFH��:��eD�*�|��N�zV�dpP�I�,(�P�xKs�Sf%y�?I��-0=�"�!��4U�=u��w闥�ܣ��/���:;��	�Q�� ƫ!���U�V���e�Ɵ
��O󉦸��:��j�AS/(-���rJd�ui�c��>��Ԣ�IK�4;��	�;��j�zu�y���Nh���<�^��s�>] �������Yޞ6��V��D,{�$�"5
4@�~���p-�z(2�G�A�6�E^7re#
���)�ِ�6̹K1�O-�Hƫ94橇�����3{Z�@��޹@{⌵��]��.�2.��p>aҐ����aO��;��~�������̨6�~L��^2�*	�I��c DB#��Nb��^��(�j�\n�5Э�,�0n�S�qw����y5dǸ�/��GP'�W�&r��k��Լ�ϪE`/Aq�0 �_�'��c�Gu��:����'��%����r������8�u�br@���ׄ��@|/k��ƗRs�����)�;N!ۃ�x<��Q/_[�7��FB�@`�!W4������Mdm�Z���5���į��Җ��7�7Y(�99�(�= ҇���)3}�����y�vˑ��:��mN�觎����QT4��N;0�p�K�e�8-�m�Wf$�"�
�Z�K]E��/)Q������鰢I�_������P�W6��*%G�����Z0�������C��~����I��X��x3��tC���^�QCN�Eu^�_q���6�{��U"�2mxW-��og��p��750������ux	����O������Lwqeh�	��NT(����|���Y%��!��1&Ǫ����rp�t��m�=��/:&�\QXvg�AC�/��;����|��':�4�#�IT�i�J���w�0���f�N2>_��h1v�]�J¶�n�9M���{+	�[�#I/��c��X��a�4��$���c� [-�N�*������)B�Vf��Wn��aAg����֩O5. Eq��J.5��O����,'8�f��A)'ZX��U�	��
uƁX�F}�>�]��R�s��2w�7`�5�������/��>�ͣm4G7N	��$��x����w�`�e-��ܮ��<V2>��8]���f�vx���p��x��'ֶ�x�Ś�8���Q�9��w���i`>��iqH�/.���p8[�jVE1"�L����.�
U�(�O�B��u�����8��=�2][gb�����Xژ!?W�^jv~̰�;v�ŏ^�z9�''��-�sb2�[�;�VT��C�Ҙ���Bƚ��yq�MXU�u�����|(���ok�������y}b�Uv�׋�r�%�v�(_��eη�4�Ӷ��C��^4𕓬7\�D���r<r�,�p��Y<&��A�VS��V���]ay��wV�k۠��SI�?�l��3��	�5^��Z"����U^%��k4�/���q����q �}a}���%�ւ�߇�E�����ռ��c��v�S�M��|ׯ���9�`z�$2ѱs��|JJ�@0���K�H8�����|��#����x�OGó߮�G���4I���{��K�gX�?��~�1�_NmA��2�d�����c<�,-�x�7Qŀh/�}����u�A�y���)�K(���U0�V�#g�۪�ͧ�"�4�Gٯ`�����T��$+;��Z`S�Pw���		ko����Ys�<L��%X��ڗ� ����H�8ןA�
�/-���6�����oD@n�������7d�Lْ�ZJ��g�8� 6o%��ퟫ��fDq@2�KD�u�Q�]!0Fqz��x�Y �͓��f��I<|lw������_=��r���d��X�%�ق�r�Y�T�"<!�2���4�Q���������5�6�?�$�z�Ď\�ٮ, ����=������ ��T��u���5Ӥ���8`�fz���|�n���������7뀦��T�Ƥ��.�
��xsi���e���XB,�{R�t��5�o[���t�%h������I�cf��Fw���J��۲1P)�>�Y�X���Y�+� �.��m8��.��k$ߵ�����}�L�)�\��}{�����Qs�����J�(���I��׼��-��Пv�Ҫ��vPP8��Bv�`�Q��j^�!9P>B�6h�B )���%6gI��Ff8n����	�Ň�rii�����s���C�}�{��m\���K��+m��.�SB��L�ڵ�[��D����n��X6l���9��nO'����J�q1��\��F��CIy|~����)���4f��*衂�[��2��r�~u�|������;�ujy����Ǵ읕���/XDD����;U�+��_��n$�S���vv���T�����X"�O��鈬o�74�E_�V3����x66D�`���N�*��e�J���+1³7�dFe�O�K���Z��H��/�Ff��6��"�
j��\�*�bI �l>���o&����w��L�b��6�z>9�����00�#^�Kdґ��n_�:�ec�����ʲ��!�T���w��Q���]R��b����e?;�m�I(�������H��)�ikU�\�<)����t6x��l^T����0�u� 2B�G�_\�u�w	E�v�FD&�"�
Ƚ�H�V~�:�h<|�7���Bg�}S�L%fe��ܤ�L�p�_:�=#��J�x�&����ZL�ߌ'���B����W� E� 3*�ﭥz�M֛XQq� D
�7�r��0E�q����UJ����Z��<;OG!F��cVY��B&��f�n,N�B�ϣ��׳.��;����澸�7Y��v;�������O
M�L�^��)[e��1$����1�ra�G�i��*�])��Ns�2���e9:���C\�����ԅ=�+G2"w9r��F yUQ����p������?8�O�Hi؞�z*�_�b��&7���R~4�9O
(�_�� �L�!�6*�h�����h�g����?�ڶ J]�f����g�LO��v��{Si��@��OU����60DI�~H��\���I�u��^c�.�XM�L�$�qm��5w|�[m�6ak׸�R�}1����_Q{��������͌��2[y��-��J���&��f%[��b�N��7��R�N&I�.xH.E5� �����~�E�c�"*�ϩ����udcB�%B�U���Z�?�Z��5�Tj��4Ns8퉹��U�m(Qy�5,:��]��\lp���p�,gC0�amo�y��[ϰq�p��
/)g+􇙔��"�J֪%�gs�K��fKU�"���K�}�#�I������u�D]J��V�e���?�D�(�W9M�Q���Jq݄��vי	������\;��3>�Ə�
�w���U�G(��u���C����ׇ�V�r��(�e������0�3�B��AeU�|�g
E'��OL��_��F���=i\�ĝ$�[�hC�u�hM��KY�ڕui����J�Tie���V{�
�u)Bu%B�"�6~�U�:��r�|���}f��y�����m��Kk
�գ��B�~۾Գ!�fdk��4=��v"����9{�+��by�F}�l��x���C��.(��ܸ�
O�1ݚ������w�g�`�?+��Ƅ�����>�����bUb��!� ���QJ���[�q�Kb��[u��Vp#c�;z������+���W�����ͬ�S��_�±�"M�C��o������*0�sw� ���j�v�-����>yMg�n$��|⃸ti��S*i\��/���`��ڵ�=�����g�d1��]�˝��xU��&�MG��|�d�>�+}�ǃ���b�ya��̴5��%�˟�FR�n;E�#�v�3}��ݚJ��Lc5?��V�@�xP`����-<� �`WQ�x�S��xw�M��sA�FV��&�x;C �*�*�V׳9���p/\)��ƨ�)��#;���q�x��v��z�K�u�8�����I�u�׌����d$����z}�i��+{�ǁ��R{E~�F�5�@,�N4��i_�ǫ�о"�u|WR�dM�`�I���`$)�B�Ճ��t�\�^p�3y"+H�9τ��4�n�E���C������Upm�ѠQ��U����ifru$-���f�Y9o�g�,OKa��`����-��L[i�c���B�=�a����3�{6� ��p����+�r??,��=wh�z�c���L�Gf+u������A����zKP�C���A��Q��!��x��f�qX�5K�<���/o�0���85#�ԝ� �����S۞����8ɚ��u�-q��1h1Y����+$�c���V����^�d�E��Ñ�.�PI�!q�gԥ^����'�V'���#m*��NWC^��[��!��#F̙�;�w�$��mf@>�����y(���H�Q�U��*���Y�*�YԮ'L�t_q�yЯ^�,�Ɖ(��/�F���P��Q��3�m�䮹�o�}K

��*�uQ��2���+L��WN�A����0e���1�٬Z��"�cZ�n
J��g�R
�����F��B�����o�����\�XM��α�e�X;/��c��@���O8�ic��P���(�B��+;�ʗ�]7�T�u@*"oG��������s�\R^���̲-�8.��-L�GeT���R
�ˋ9Vs������Ŀ���:�d!�kJ�u��q�E0���.[�Y/��^/}��󮘾�R�ܓ��P�V�~u�?ö4��5A*���Ɍ�����<��Uhj�Y�;���*���)�c�X��1�U�����Z1g7�p��#�1��U:�C%�N��5�(�cȵ��񦰈?�ӭ�w�����������䵔.��p�h<��"(/u�(}��
G�g��T�[�I��H_��7�A��WlK���O��,*Vh_�Pih3}�7_�LM�t�hZĽo��)�-gI`��?O��W�Xf������^V���B����S��j�y,<5}�W ����'�Z��+�ψ@]KK��Ci�ۑZњM��/��*L�r�>���M S3�G����	����`d
��P�O�$��L� ���4�Ó�3�I@�.Α-S�2���i艶ͥ���F�T^Y�MtOL�+T#~�	�W�����!�P�;_�7��~���]��X���5p�"�>"��<�+����i �L_ظ�Bݬ2�v��ٳ�[�ޅ$�-��̬7���5X�~$�s�ʓ�C�����y���A�Fn�e��2����,JI6���.�
�t�Ø_�����0�5Zd��θ�����`����<�X�<�
PN�i�p_?�WK��~x��?�qO��7�P� �������oV��'��=�Ӯ��_����gDY��%�|��#��c� :sv�5���0�e7��F�%�|��kZ�)ʘ\�j}I;z��RvM� �eQi9�==�Ǌ�Zym�ˊ��g1gq�y@�3��c��t#�Ky� ��oٗ=0Mq�w�MY���ݩ��L9�"D�m�>3����[�~�8�,�M���^��Be=�	��'�~�8��F�D����}U��G�_�0>�(CJ�j�{�Ǯ��$��H�_)�V|����yo�,���ԩ�0fT��`J��w�	w�¹��u� ]:Q�뙏�ޛ�0�w��X�����|��k��	��%m�@��)�W��rnU�ӷ��¸��m��]���ev�8/��2��«ǰ����S�pK�
�q����f��>����%H!-G!�����/>��ok�M�xt�՝_�~K$j=(�PK   !l�Y�_���  �     jsons/user_defined.json��]o�6����kS��7s���M�8
lA!QT*��<�^��;��-M�n�+Y"�C�}��/��q�l������M�l����Mӵ���4��ٕC�Mv�Ǘ�?W�����������[>{�|g�R��[����>�l��o�v�ճ�OM{����c��>�ٶ��y��Uf\�A��x[[µ�t�.,����*�2��߸�Yo�Ѿ��8�_W�5�@���D����"�Ђ�V
���=�k\�N�lYִ�N�JE������)WزpB8��顸��;|�)�
/W]�>y|�n�˶/Y�{X4���x��V��l.���<��>��0��oBL)ߵ�_;|���Zn{���m�ݦ��iVx�I@,�0����h6������9ѫ��C�s�=��!��	�y^��W�_�Q<�b�K���}��.:��J_�(]t5���d:��e@���d:D�*��13R�d�E�����&��S�t�^$���oQ��0�Y�<6�!�+L���~��jF�Za�g櫫8?-��U�&Ϟ��M<@�[�#������5eH�=�{��{� �z�097F��+���G��W��'>����=@�`1�������@�`D:��B�q�Z�t��/[���4~���cf��̀��Kj��o(b;����8�����	��)��h� ��
�@��6����x�P��Ǐ,x�K\�U���H�E7GX�'SH���iz`5���+yT�ݸ���
��M����껵��X�`�=��ַ������}[�9��)P6���vv�Eάh����};[�v��A���m�<�6��T��W�Т.�H��P*� J�"��)uQ��FDآ���rRV�jg$2��k����8T�ȜS&~�r�2W��ޜ��=j�H�r{yd�rh��M�z�n$W��[��'T.l�g����	���Ҥ�/��[��<�~��������E��:7��7՞.R��9�ˉ Պ���A��R^�r8�(�s�2@]Y�U�d#4���l�����wf�=b�lw{����Ea�H��_U�"J�-X��hB4����ķ"P�c��W+�-<Ȋ��''��JZk*M%�����1S��Q��''�=��>xr9eZ����[4 �e�9ڻʥ6�T�ւ��������S�O��tR��E�mH�@���R��t��/PK
   !l�Y^!H��  �a                   cirkitFile.jsonPK
   lg�YG���F"  A"  /               images/07631829-c1ba-46e6-b58f-b7cc9d810cbd.pngPK
   �f�Y�7}b  ]  /             �.  images/9bbf0d51-8956-46f1-ad90-c6ca9bac44cc.pngPK
   lg�Y�{�" %# /             SG  images/b7ab4f1c-086a-49aa-bc93-bd307c85ad93.pngPK
   Th�Y����  (  /             �_ images/c33d050f-98d7-424b-970e-349228d04709.pngPK
   Th�Y��:$  �  /             | images/f2ef8506-1b6f-4eaa-8cf6-e59ae15d09b8.pngPK
   �f�Y8�w���  ��  /             �� images/fd1e7351-dbfe-4fec-861d-4a74217661c3.pngPK
   !l�Y�_���  �               �g jsons/user_defined.jsonPK      �  �l   